module wen_in_1_reg_value (
    input [28:0] I,
    output [0:0] O
);
assign O = I[28];
endmodule

module wen_in_1_reg_sel (
    input [28:0] I,
    output [0:0] O
);
assign O = I[27];
endmodule

module wen_in_0_reg_value (
    input [28:0] I,
    output [0:0] O
);
assign O = I[26];
endmodule

module wen_in_0_reg_sel (
    input [28:0] I,
    output [0:0] O
);
assign O = I[25];
endmodule

module tile_en (
    input [28:0] I,
    output [0:0] O
);
assign O = I[24];
endmodule

module strg_ub_tb_only_tb_write_addr_gen_1_strides_5 (
    input [28:0] I,
    output [3:0] O
);
assign O = I[23:20];
endmodule

module strg_ub_tb_only_tb_write_addr_gen_1_strides_4 (
    input [28:0] I,
    output [3:0] O
);
assign O = I[19:16];
endmodule

module strg_ub_tb_only_tb_write_addr_gen_1_strides_3 (
    input [28:0] I,
    output [3:0] O
);
assign O = I[15:12];
endmodule

module strg_ub_tb_only_tb_write_addr_gen_1_strides_2 (
    input [28:0] I,
    output [3:0] O
);
assign O = I[11:8];
endmodule

module strg_ub_tb_only_tb_write_addr_gen_1_strides_1 (
    input [28:0] I,
    output [3:0] O
);
assign O = I[7:4];
endmodule

module strg_ub_tb_only_tb_write_addr_gen_1_strides_0 (
    input [28:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module strg_ub_tb_only_tb_write_addr_gen_1_starting_addr (
    input [31:0] I,
    output [3:0] O
);
assign O = I[31:28];
endmodule

module strg_ub_tb_only_tb_write_addr_gen_0_strides_5 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[27:24];
endmodule

module strg_ub_tb_only_tb_write_addr_gen_0_strides_4 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[23:20];
endmodule

module strg_ub_tb_only_tb_write_addr_gen_0_strides_3 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[19:16];
endmodule

module strg_ub_tb_only_tb_write_addr_gen_0_strides_2 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[15:12];
endmodule

module strg_ub_tb_only_tb_write_addr_gen_0_strides_1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[11:8];
endmodule

module strg_ub_tb_only_tb_write_addr_gen_0_strides_0 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[7:4];
endmodule

module strg_ub_tb_only_tb_write_addr_gen_0_starting_addr (
    input [31:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr (
    input [16:0] I,
    output [15:0] O
);
assign O = I[16:1];
endmodule

module strg_ub_tb_only_tb_read_sched_gen_1_enable (
    input [16:0] I,
    output [0:0] O
);
assign O = I[0];
endmodule

module strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr (
    input [24:0] I,
    output [15:0] O
);
assign O = I[24:9];
endmodule

module strg_ub_tb_only_tb_read_sched_gen_0_enable (
    input [24:0] I,
    output [0:0] O
);
assign O = I[8];
endmodule

module strg_ub_tb_only_tb_read_addr_gen_1_strides_5 (
    input [24:0] I,
    output [3:0] O
);
assign O = I[7:4];
endmodule

module strg_ub_tb_only_tb_read_addr_gen_1_strides_4 (
    input [24:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module strg_ub_tb_only_tb_read_addr_gen_1_strides_3 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[31:28];
endmodule

module strg_ub_tb_only_tb_read_addr_gen_1_strides_2 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[27:24];
endmodule

module strg_ub_tb_only_tb_read_addr_gen_1_strides_1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[23:20];
endmodule

module strg_ub_tb_only_tb_read_addr_gen_1_strides_0 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[19:16];
endmodule

module strg_ub_tb_only_tb_read_addr_gen_1_starting_addr (
    input [31:0] I,
    output [3:0] O
);
assign O = I[15:12];
endmodule

module strg_ub_tb_only_tb_read_addr_gen_0_strides_5 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[11:8];
endmodule

module strg_ub_tb_only_tb_read_addr_gen_0_strides_4 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[7:4];
endmodule

module strg_ub_tb_only_tb_read_addr_gen_0_strides_3 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module strg_ub_tb_only_tb_read_addr_gen_0_strides_2 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[31:28];
endmodule

module strg_ub_tb_only_tb_read_addr_gen_0_strides_1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[27:24];
endmodule

module strg_ub_tb_only_tb_read_addr_gen_0_strides_0 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[23:20];
endmodule

module strg_ub_tb_only_tb_read_addr_gen_0_starting_addr (
    input [31:0] I,
    output [3:0] O
);
assign O = I[19:16];
endmodule

module strg_ub_tb_only_loops_buf2out_read_1_ranges_5 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_tb_only_loops_buf2out_read_1_ranges_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_tb_only_loops_buf2out_read_1_ranges_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_tb_only_loops_buf2out_read_1_ranges_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_tb_only_loops_buf2out_read_1_ranges_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_tb_only_loops_buf2out_read_1_ranges_0 (
    input [19:0] I,
    output [15:0] O
);
assign O = I[19:4];
endmodule

module strg_ub_tb_only_loops_buf2out_read_1_dimensionality (
    input [19:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module strg_ub_tb_only_loops_buf2out_read_0_ranges_5 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_tb_only_loops_buf2out_read_0_ranges_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_tb_only_loops_buf2out_read_0_ranges_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_tb_only_loops_buf2out_read_0_ranges_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_tb_only_loops_buf2out_read_0_ranges_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_tb_only_loops_buf2out_read_0_ranges_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_tb_only_loops_buf2out_read_0_dimensionality (
    input [19:0] I,
    output [3:0] O
);
assign O = I[19:16];
endmodule

module strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5 (
    input [19:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_sram_tb_shared_output_sched_gen_1_enable (
    input [16:0] I,
    output [0:0] O
);
assign O = I[16];
endmodule

module strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5 (
    input [16:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_sram_tb_shared_output_sched_gen_0_enable (
    input [16:0] I,
    output [0:0] O
);
assign O = I[16];
endmodule

module strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5 (
    input [16:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0 (
    input [19:0] I,
    output [15:0] O
);
assign O = I[19:4];
endmodule

module strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality (
    input [19:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality (
    input [30:0] I,
    output [3:0] O
);
assign O = I[30:27];
endmodule

module strg_ub_sram_only_output_addr_gen_1_strides_5 (
    input [30:0] I,
    output [8:0] O
);
assign O = I[26:18];
endmodule

module strg_ub_sram_only_output_addr_gen_1_strides_4 (
    input [30:0] I,
    output [8:0] O
);
assign O = I[17:9];
endmodule

module strg_ub_sram_only_output_addr_gen_1_strides_3 (
    input [30:0] I,
    output [8:0] O
);
assign O = I[8:0];
endmodule

module strg_ub_sram_only_output_addr_gen_1_strides_2 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[26:18];
endmodule

module strg_ub_sram_only_output_addr_gen_1_strides_1 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[17:9];
endmodule

module strg_ub_sram_only_output_addr_gen_1_strides_0 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[8:0];
endmodule

module strg_ub_sram_only_output_addr_gen_1_starting_addr (
    input [26:0] I,
    output [8:0] O
);
assign O = I[26:18];
endmodule

module strg_ub_sram_only_output_addr_gen_0_strides_5 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[17:9];
endmodule

module strg_ub_sram_only_output_addr_gen_0_strides_4 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[8:0];
endmodule

module strg_ub_sram_only_output_addr_gen_0_strides_3 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[26:18];
endmodule

module strg_ub_sram_only_output_addr_gen_0_strides_2 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[17:9];
endmodule

module strg_ub_sram_only_output_addr_gen_0_strides_1 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[8:0];
endmodule

module strg_ub_sram_only_output_addr_gen_0_strides_0 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[26:18];
endmodule

module strg_ub_sram_only_output_addr_gen_0_starting_addr (
    input [26:0] I,
    output [8:0] O
);
assign O = I[17:9];
endmodule

module strg_ub_sram_only_input_addr_gen_1_strides_5 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[8:0];
endmodule

module strg_ub_sram_only_input_addr_gen_1_strides_4 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[26:18];
endmodule

module strg_ub_sram_only_input_addr_gen_1_strides_3 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[17:9];
endmodule

module strg_ub_sram_only_input_addr_gen_1_strides_2 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[8:0];
endmodule

module strg_ub_sram_only_input_addr_gen_1_strides_1 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[26:18];
endmodule

module strg_ub_sram_only_input_addr_gen_1_strides_0 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[17:9];
endmodule

module strg_ub_sram_only_input_addr_gen_1_starting_addr (
    input [26:0] I,
    output [8:0] O
);
assign O = I[8:0];
endmodule

module strg_ub_sram_only_input_addr_gen_0_strides_5 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[26:18];
endmodule

module strg_ub_sram_only_input_addr_gen_0_strides_4 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[17:9];
endmodule

module strg_ub_sram_only_input_addr_gen_0_strides_3 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[8:0];
endmodule

module strg_ub_sram_only_input_addr_gen_0_strides_2 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[26:18];
endmodule

module strg_ub_sram_only_input_addr_gen_0_strides_1 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[17:9];
endmodule

module strg_ub_sram_only_input_addr_gen_0_strides_0 (
    input [26:0] I,
    output [8:0] O
);
assign O = I[8:0];
endmodule

module strg_ub_sram_only_input_addr_gen_0_starting_addr (
    input [24:0] I,
    output [8:0] O
);
assign O = I[24:16];
endmodule

module strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5 (
    input [24:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0 (
    input [19:0] I,
    output [15:0] O
);
assign O = I[19:4];
endmodule

module strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality (
    input [19:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality (
    input [19:0] I,
    output [3:0] O
);
assign O = I[19:16];
endmodule

module strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5 (
    input [19:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_sram_shared_agg_read_sched_gen_1_enable (
    input [16:0] I,
    output [0:0] O
);
assign O = I[16];
endmodule

module strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5 (
    input [16:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_sram_shared_agg_read_sched_gen_0_enable (
    input [16:0] I,
    output [0:0] O
);
assign O = I[16];
endmodule

module strg_ub_agg_only_loops_in2buf_1_ranges_5 (
    input [16:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_only_loops_in2buf_1_ranges_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_agg_only_loops_in2buf_1_ranges_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_only_loops_in2buf_1_ranges_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_agg_only_loops_in2buf_1_ranges_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_only_loops_in2buf_1_ranges_0 (
    input [19:0] I,
    output [15:0] O
);
assign O = I[19:4];
endmodule

module strg_ub_agg_only_loops_in2buf_1_dimensionality (
    input [19:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module strg_ub_agg_only_loops_in2buf_0_ranges_5 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_agg_only_loops_in2buf_0_ranges_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_only_loops_in2buf_0_ranges_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_agg_only_loops_in2buf_0_ranges_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_only_loops_in2buf_0_ranges_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_agg_only_loops_in2buf_0_ranges_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_only_loops_in2buf_0_dimensionality (
    input [19:0] I,
    output [3:0] O
);
assign O = I[19:16];
endmodule

module strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5 (
    input [19:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_only_agg_write_sched_gen_1_enable (
    input [16:0] I,
    output [0:0] O
);
assign O = I[16];
endmodule

module strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5 (
    input [16:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module strg_ub_agg_only_agg_write_sched_gen_0_enable (
    input [16:0] I,
    output [0:0] O
);
assign O = I[16];
endmodule

module strg_ub_agg_only_agg_write_addr_gen_1_strides_5 (
    input [16:0] I,
    output [3:0] O
);
assign O = I[15:12];
endmodule

module strg_ub_agg_only_agg_write_addr_gen_1_strides_4 (
    input [16:0] I,
    output [3:0] O
);
assign O = I[11:8];
endmodule

module strg_ub_agg_only_agg_write_addr_gen_1_strides_3 (
    input [16:0] I,
    output [3:0] O
);
assign O = I[7:4];
endmodule

module strg_ub_agg_only_agg_write_addr_gen_1_strides_2 (
    input [16:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module strg_ub_agg_only_agg_write_addr_gen_1_strides_1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[31:28];
endmodule

module strg_ub_agg_only_agg_write_addr_gen_1_strides_0 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[27:24];
endmodule

module strg_ub_agg_only_agg_write_addr_gen_1_starting_addr (
    input [31:0] I,
    output [3:0] O
);
assign O = I[23:20];
endmodule

module strg_ub_agg_only_agg_write_addr_gen_0_strides_5 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[19:16];
endmodule

module strg_ub_agg_only_agg_write_addr_gen_0_strides_4 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[15:12];
endmodule

module strg_ub_agg_only_agg_write_addr_gen_0_strides_3 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[11:8];
endmodule

module strg_ub_agg_only_agg_write_addr_gen_0_strides_2 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[7:4];
endmodule

module strg_ub_agg_only_agg_write_addr_gen_0_strides_1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module strg_ub_agg_only_agg_write_addr_gen_0_strides_0 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[31:28];
endmodule

module strg_ub_agg_only_agg_write_addr_gen_0_starting_addr (
    input [31:0] I,
    output [3:0] O
);
assign O = I[27:24];
endmodule

module strg_ub_agg_only_agg_read_addr_gen_1_strides_5 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[23:20];
endmodule

module strg_ub_agg_only_agg_read_addr_gen_1_strides_4 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[19:16];
endmodule

module strg_ub_agg_only_agg_read_addr_gen_1_strides_3 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[15:12];
endmodule

module strg_ub_agg_only_agg_read_addr_gen_1_strides_2 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[11:8];
endmodule

module strg_ub_agg_only_agg_read_addr_gen_1_strides_1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[7:4];
endmodule

module strg_ub_agg_only_agg_read_addr_gen_1_strides_0 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module strg_ub_agg_only_agg_read_addr_gen_1_starting_addr (
    input [31:0] I,
    output [3:0] O
);
assign O = I[31:28];
endmodule

module strg_ub_agg_only_agg_read_addr_gen_0_strides_5 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[27:24];
endmodule

module strg_ub_agg_only_agg_read_addr_gen_0_strides_4 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[23:20];
endmodule

module strg_ub_agg_only_agg_read_addr_gen_0_strides_3 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[19:16];
endmodule

module strg_ub_agg_only_agg_read_addr_gen_0_strides_2 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[15:12];
endmodule

module strg_ub_agg_only_agg_read_addr_gen_0_strides_1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[11:8];
endmodule

module strg_ub_agg_only_agg_read_addr_gen_0_strides_0 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[7:4];
endmodule

module strg_ub_agg_only_agg_read_addr_gen_0_starting_addr (
    input [31:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module stencil_valid_sched_gen_sched_addr_gen_strides_5 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module stencil_valid_sched_gen_sched_addr_gen_strides_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module stencil_valid_sched_gen_sched_addr_gen_strides_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module stencil_valid_sched_gen_sched_addr_gen_strides_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module stencil_valid_sched_gen_sched_addr_gen_strides_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module stencil_valid_sched_gen_sched_addr_gen_strides_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module stencil_valid_sched_gen_sched_addr_gen_starting_addr (
    input [22:0] I,
    output [15:0] O
);
assign O = I[22:7];
endmodule

module stencil_valid_sched_gen_enable (
    input [22:0] I,
    output [0:0] O
);
assign O = I[6];
endmodule

module ren_in_1_reg_value (
    input [22:0] I,
    output [0:0] O
);
assign O = I[5];
endmodule

module ren_in_1_reg_sel (
    input [22:0] I,
    output [0:0] O
);
assign O = I[4];
endmodule

module ren_in_0_reg_value (
    input [22:0] I,
    output [0:0] O
);
assign O = I[3];
endmodule

module ren_in_0_reg_sel (
    input [22:0] I,
    output [0:0] O
);
assign O = I[2];
endmodule

module mode (
    input [22:0] I,
    output [1:0] O
);
assign O = I[1:0];
endmodule

module mantle_wire__typeBitIn8 (
    output [7:0] in,
    input [7:0] out
);
assign in = out;
endmodule

module mantle_wire__typeBitIn7 (
    output [6:0] in,
    input [6:0] out
);
assign in = out;
endmodule

module mantle_wire__typeBitIn4 (
    output [3:0] in,
    input [3:0] out
);
assign in = out;
endmodule

module mantle_wire__typeBitIn32 (
    output [31:0] in,
    input [31:0] out
);
assign in = out;
endmodule

module mantle_wire__typeBitIn2 (
    output [1:0] in,
    input [1:0] out
);
assign in = out;
endmodule

module mantle_wire__typeBitIn16 (
    output [15:0] in,
    input [15:0] out
);
assign in = out;
endmodule

module mantle_wire__typeBit9 (
    input [8:0] in,
    output [8:0] out
);
assign out = in;
endmodule

module mantle_wire__typeBit8 (
    input [7:0] in,
    output [7:0] out
);
assign out = in;
endmodule

module mantle_wire__typeBit5 (
    input [4:0] in,
    output [4:0] out
);
assign out = in;
endmodule

module mantle_wire__typeBit4 (
    input [3:0] in,
    output [3:0] out
);
assign out = in;
endmodule

module mantle_wire__typeBit32 (
    input [31:0] in,
    output [31:0] out
);
assign out = in;
endmodule

module mantle_wire__typeBit31 (
    input [30:0] in,
    output [30:0] out
);
assign out = in;
endmodule

module mantle_wire__typeBit30 (
    input [29:0] in,
    output [29:0] out
);
assign out = in;
endmodule

module mantle_wire__typeBit29 (
    input [28:0] in,
    output [28:0] out
);
assign out = in;
endmodule

module mantle_wire__typeBit28 (
    input [27:0] in,
    output [27:0] out
);
assign out = in;
endmodule

module mantle_wire__typeBit27 (
    input [26:0] in,
    output [26:0] out
);
assign out = in;
endmodule

module mantle_wire__typeBit25 (
    input [24:0] in,
    output [24:0] out
);
assign out = in;
endmodule

module mantle_wire__typeBit23 (
    input [22:0] in,
    output [22:0] out
);
assign out = in;
endmodule

module mantle_wire__typeBit20 (
    input [19:0] in,
    output [19:0] out
);
assign out = in;
endmodule

module mantle_wire__typeBit18 (
    input [17:0] in,
    output [17:0] out
);
assign out = in;
endmodule

module mantle_wire__typeBit17 (
    input [16:0] in,
    output [16:0] out
);
assign out = in;
endmodule

module mantle_wire__typeBit16 (
    input [15:0] in,
    output [15:0] out
);
assign out = in;
endmodule

module regCE_arst #(
    parameter width = 1,
    parameter init = 1
) (
    input [width-1:0] in,
    input ce,
    output [width-1:0] out,
    input clk,
    input arst
);
  reg [width-1:0] value;
  always @(posedge clk, posedge arst) begin
    if (arst) begin
      value <= init;
    end
    else if (ce) begin
      value <= in;
    end
  end
  assign out = value;
endmodule

module regCE #(
    parameter width = 1
) (
    input [width-1:0] in,
    input ce,
    output [width-1:0] out,
    input clk
);
  reg [width-1:0] value;
  always @(posedge clk) begin
    if (ce) begin
      value <= in;
    end
  end
  assign out = value;
endmodule

module loops_stencil_valid_ranges_5 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module loops_stencil_valid_ranges_4 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module loops_stencil_valid_ranges_3 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module loops_stencil_valid_ranges_2 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module loops_stencil_valid_ranges_1 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[31:16];
endmodule

module loops_stencil_valid_ranges_0 (
    input [31:0] I,
    output [15:0] O
);
assign O = I[15:0];
endmodule

module loops_stencil_valid_dimensionality (
    input [22:0] I,
    output [3:0] O
);
assign O = I[22:19];
endmodule

module io_core (
    input [15:0] glb2io_16,
    input [0:0] glb2io_1,
    output [15:0] io2glb_16,
    output [0:0] io2glb_1,
    input [15:0] f2io_16,
    input [0:0] f2io_1,
    output [15:0] io2f_16,
    output [0:0] io2f_1
);
assign io2glb_16 = f2io_16;
assign io2glb_1 = f2io_1;
assign io2f_16 = glb2io_16;
assign io2f_1 = glb2io_1;
endmodule

module inst_1 (
    input [31:0] I,
    output [31:0] O
);
assign O = I;
endmodule

module inst_0 (
    input [31:0] I,
    output [31:0] O
);
assign O = I;
endmodule

module flush_reg_value (
    input [22:0] I,
    output [0:0] O
);
assign O = I[18];
endmodule

module flush_reg_sel (
    input [22:0] I,
    output [0:0] O
);
assign O = I[17];
endmodule

module fifo_ctrl_fifo_depth (
    input [22:0] I,
    output [15:0] O
);
assign O = I[16:1];
endmodule

module coreir_xor #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output [width-1:0] out
);
  assign out = in0 ^ in1;
endmodule

module coreir_wrap (
    input in,
    output out
);
  assign out = in;
endmodule

module coreir_ult #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output out
);
  assign out = in0 < in1;
endmodule

module coreir_ule #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output out
);
  assign out = in0 <= in1;
endmodule

module coreir_uge #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output out
);
  assign out = in0 >= in1;
endmodule

module coreir_slt #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output out
);
  assign out = $signed(in0) < $signed(in1);
endmodule

module coreir_slice #(
    parameter hi = 1,
    parameter lo = 0,
    parameter width = 1
) (
    input [width-1:0] in,
    output [hi-lo-1:0] out
);
  assign out = in[hi-1:lo];
endmodule

module coreir_sle #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output out
);
  assign out = $signed(in0) <= $signed(in1);
endmodule

module coreir_sge #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output out
);
  assign out = $signed(in0) >= $signed(in1);
endmodule

module coreir_reg #(
    parameter width = 1,
    parameter clk_posedge = 1,
    parameter init = 1
) (
    input clk,
    input [width-1:0] in,
    output [width-1:0] out
);
  reg [width-1:0] outReg=init;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk) begin
    outReg <= in;
  end
  assign out = outReg;
endmodule

module coreir_orr #(
    parameter width = 1
) (
    input [width-1:0] in,
    output out
);
  assign out = |in;
endmodule

module coreir_or #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output [width-1:0] out
);
  assign out = in0 | in1;
endmodule

module coreir_not #(
    parameter width = 1
) (
    input [width-1:0] in,
    output [width-1:0] out
);
  assign out = ~in;
endmodule

module coreir_neg #(
    parameter width = 1
) (
    input [width-1:0] in,
    output [width-1:0] out
);
  assign out = -in;
endmodule

module coreir_mux #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    input sel,
    output [width-1:0] out
);
  assign out = sel ? in1 : in0;
endmodule

module coreir_mul #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output [width-1:0] out
);
  assign out = in0 * in1;
endmodule

module coreir_lshr #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output [width-1:0] out
);
  assign out = in0 >> in1;
endmodule

module coreir_eq #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output out
);
  assign out = in0 == in1;
endmodule

module coreir_const #(
    parameter width = 1,
    parameter value = 1
) (
    output [width-1:0] out
);
  assign out = value;
endmodule

module coreir_ashr #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output [width-1:0] out
);
  assign out = $signed(in0) >>> in1;
endmodule

module coreir_and #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output [width-1:0] out
);
  assign out = in0 & in1;
endmodule

module coreir_add #(
    parameter width = 1
) (
    input [width-1:0] in0,
    input [width-1:0] in1,
    output [width-1:0] out
);
  assign out = in0 + in1;
endmodule

module corebit_xor (
    input in0,
    input in1,
    output out
);
  assign out = in0 ^ in1;
endmodule

module corebit_term (
    input in
);

endmodule

module corebit_or (
    input in0,
    input in1,
    output out
);
  assign out = in0 | in1;
endmodule

module corebit_not (
    input in,
    output out
);
  assign out = ~in;
endmodule

module corebit_const #(
    parameter value = 1
) (
    output out
);
  assign out = value;
endmodule

module corebit_and (
    input in0,
    input in1,
    output out
);
  assign out = in0 & in1;
endmodule

module commonlib_muxn__N2__width32 (
    input [31:0] in_data_0,
    input [31:0] in_data_1,
    input [0:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
coreir_mux #(
    .width(32)
) _join (
    .in0(in_data_0),
    .in1(in_data_1),
    .sel(in_sel[0]),
    .out(_join_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N4__width32 (
    input [31:0] in_data_0,
    input [31:0] in_data_1,
    input [31:0] in_data_2,
    input [31:0] in_data_3,
    input [1:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
wire [31:0] muxN_0_out;
wire [31:0] muxN_1_out;
wire [0:0] sel_slice0_out;
wire [0:0] sel_slice1_out;
coreir_mux #(
    .width(32)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[1]),
    .out(_join_out)
);
commonlib_muxn__N2__width32 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N2__width32 muxN_1 (
    .in_data_0(in_data_2),
    .in_data_1(in_data_3),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(1),
    .lo(0),
    .width(2)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(1),
    .lo(0),
    .width(2)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N8__width32 (
    input [31:0] in_data_0,
    input [31:0] in_data_1,
    input [31:0] in_data_2,
    input [31:0] in_data_3,
    input [31:0] in_data_4,
    input [31:0] in_data_5,
    input [31:0] in_data_6,
    input [31:0] in_data_7,
    input [2:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
wire [31:0] muxN_0_out;
wire [31:0] muxN_1_out;
wire [1:0] sel_slice0_out;
wire [1:0] sel_slice1_out;
coreir_mux #(
    .width(32)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[2]),
    .out(_join_out)
);
commonlib_muxn__N4__width32 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_2(in_data_2),
    .in_data_3(in_data_3),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N4__width32 muxN_1 (
    .in_data_0(in_data_4),
    .in_data_1(in_data_5),
    .in_data_2(in_data_6),
    .in_data_3(in_data_7),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(2),
    .lo(0),
    .width(3)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(2),
    .lo(0),
    .width(3)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N2__width16 (
    input [15:0] in_data_0,
    input [15:0] in_data_1,
    input [0:0] in_sel,
    output [15:0] out
);
wire [15:0] _join_out;
coreir_mux #(
    .width(16)
) _join (
    .in0(in_data_0),
    .in1(in_data_1),
    .sel(in_sel[0]),
    .out(_join_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N4__width16 (
    input [15:0] in_data_0,
    input [15:0] in_data_1,
    input [15:0] in_data_2,
    input [15:0] in_data_3,
    input [1:0] in_sel,
    output [15:0] out
);
wire [15:0] _join_out;
wire [15:0] muxN_0_out;
wire [15:0] muxN_1_out;
wire [0:0] sel_slice0_out;
wire [0:0] sel_slice1_out;
coreir_mux #(
    .width(16)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[1]),
    .out(_join_out)
);
commonlib_muxn__N2__width16 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N2__width16 muxN_1 (
    .in_data_0(in_data_2),
    .in_data_1(in_data_3),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(1),
    .lo(0),
    .width(2)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(1),
    .lo(0),
    .width(2)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N8__width16 (
    input [15:0] in_data_0,
    input [15:0] in_data_1,
    input [15:0] in_data_2,
    input [15:0] in_data_3,
    input [15:0] in_data_4,
    input [15:0] in_data_5,
    input [15:0] in_data_6,
    input [15:0] in_data_7,
    input [2:0] in_sel,
    output [15:0] out
);
wire [15:0] _join_out;
wire [15:0] muxN_0_out;
wire [15:0] muxN_1_out;
wire [1:0] sel_slice0_out;
wire [1:0] sel_slice1_out;
coreir_mux #(
    .width(16)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[2]),
    .out(_join_out)
);
commonlib_muxn__N4__width16 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_2(in_data_2),
    .in_data_3(in_data_3),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N4__width16 muxN_1 (
    .in_data_0(in_data_4),
    .in_data_1(in_data_5),
    .in_data_2(in_data_6),
    .in_data_3(in_data_7),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(2),
    .lo(0),
    .width(3)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(2),
    .lo(0),
    .width(3)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N2__width1 (
    input [0:0] in_data_0,
    input [0:0] in_data_1,
    input [0:0] in_sel,
    output [0:0] out
);
wire [0:0] _join_out;
coreir_mux #(
    .width(1)
) _join (
    .in0(in_data_0),
    .in1(in_data_1),
    .sel(in_sel[0]),
    .out(_join_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N4__width1 (
    input [0:0] in_data_0,
    input [0:0] in_data_1,
    input [0:0] in_data_2,
    input [0:0] in_data_3,
    input [1:0] in_sel,
    output [0:0] out
);
wire [0:0] _join_out;
wire [0:0] muxN_0_out;
wire [0:0] muxN_1_out;
wire [0:0] sel_slice0_out;
wire [0:0] sel_slice1_out;
coreir_mux #(
    .width(1)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[1]),
    .out(_join_out)
);
commonlib_muxn__N2__width1 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N2__width1 muxN_1 (
    .in_data_0(in_data_2),
    .in_data_1(in_data_3),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(1),
    .lo(0),
    .width(2)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(1),
    .lo(0),
    .width(2)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N8__width1 (
    input [0:0] in_data_0,
    input [0:0] in_data_1,
    input [0:0] in_data_2,
    input [0:0] in_data_3,
    input [0:0] in_data_4,
    input [0:0] in_data_5,
    input [0:0] in_data_6,
    input [0:0] in_data_7,
    input [2:0] in_sel,
    output [0:0] out
);
wire [0:0] _join_out;
wire [0:0] muxN_0_out;
wire [0:0] muxN_1_out;
wire [1:0] sel_slice0_out;
wire [1:0] sel_slice1_out;
coreir_mux #(
    .width(1)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[2]),
    .out(_join_out)
);
commonlib_muxn__N4__width1 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_2(in_data_2),
    .in_data_3(in_data_3),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N4__width1 muxN_1 (
    .in_data_0(in_data_4),
    .in_data_1(in_data_5),
    .in_data_2(in_data_6),
    .in_data_3(in_data_7),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(2),
    .lo(0),
    .width(3)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(2),
    .lo(0),
    .width(3)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N1__width32 (
    input [31:0] in_data_0,
    input [0:0] in_sel,
    output [31:0] out
);
corebit_term term_sel (
    .in(in_sel[0])
);
assign out = in_data_0;
endmodule

module commonlib_muxn__N9__width32 (
    input [31:0] in_data_0,
    input [31:0] in_data_1,
    input [31:0] in_data_2,
    input [31:0] in_data_3,
    input [31:0] in_data_4,
    input [31:0] in_data_5,
    input [31:0] in_data_6,
    input [31:0] in_data_7,
    input [31:0] in_data_8,
    input [3:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
wire [31:0] muxN_0_out;
wire [31:0] muxN_1_out;
wire [2:0] sel_slice0_out;
wire [0:0] sel_slice1_out;
coreir_mux #(
    .width(32)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[3]),
    .out(_join_out)
);
commonlib_muxn__N8__width32 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_2(in_data_2),
    .in_data_3(in_data_3),
    .in_data_4(in_data_4),
    .in_data_5(in_data_5),
    .in_data_6(in_data_6),
    .in_data_7(in_data_7),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N1__width32 muxN_1 (
    .in_data_0(in_data_8),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(3),
    .lo(0),
    .width(4)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(1),
    .lo(0),
    .width(4)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N3__width32 (
    input [31:0] in_data_0,
    input [31:0] in_data_1,
    input [31:0] in_data_2,
    input [1:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
wire [31:0] muxN_0_out;
wire [31:0] muxN_1_out;
wire [0:0] sel_slice0_out;
wire [0:0] sel_slice1_out;
coreir_mux #(
    .width(32)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[1]),
    .out(_join_out)
);
commonlib_muxn__N2__width32 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N1__width32 muxN_1 (
    .in_data_0(in_data_2),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(1),
    .lo(0),
    .width(2)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(1),
    .lo(0),
    .width(2)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N1__width16 (
    input [15:0] in_data_0,
    input [0:0] in_sel,
    output [15:0] out
);
corebit_term term_sel (
    .in(in_sel[0])
);
assign out = in_data_0;
endmodule

module commonlib_muxn__N5__width16 (
    input [15:0] in_data_0,
    input [15:0] in_data_1,
    input [15:0] in_data_2,
    input [15:0] in_data_3,
    input [15:0] in_data_4,
    input [2:0] in_sel,
    output [15:0] out
);
wire [15:0] _join_out;
wire [15:0] muxN_0_out;
wire [15:0] muxN_1_out;
wire [1:0] sel_slice0_out;
wire [0:0] sel_slice1_out;
coreir_mux #(
    .width(16)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[2]),
    .out(_join_out)
);
commonlib_muxn__N4__width16 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_2(in_data_2),
    .in_data_3(in_data_3),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N1__width16 muxN_1 (
    .in_data_0(in_data_4),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(2),
    .lo(0),
    .width(3)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(1),
    .lo(0),
    .width(3)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N1__width1 (
    input [0:0] in_data_0,
    input [0:0] in_sel,
    output [0:0] out
);
corebit_term term_sel (
    .in(in_sel[0])
);
assign out = in_data_0;
endmodule

module commonlib_muxn__N9__width1 (
    input [0:0] in_data_0,
    input [0:0] in_data_1,
    input [0:0] in_data_2,
    input [0:0] in_data_3,
    input [0:0] in_data_4,
    input [0:0] in_data_5,
    input [0:0] in_data_6,
    input [0:0] in_data_7,
    input [0:0] in_data_8,
    input [3:0] in_sel,
    output [0:0] out
);
wire [0:0] _join_out;
wire [0:0] muxN_0_out;
wire [0:0] muxN_1_out;
wire [2:0] sel_slice0_out;
wire [0:0] sel_slice1_out;
coreir_mux #(
    .width(1)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[3]),
    .out(_join_out)
);
commonlib_muxn__N8__width1 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_2(in_data_2),
    .in_data_3(in_data_3),
    .in_data_4(in_data_4),
    .in_data_5(in_data_5),
    .in_data_6(in_data_6),
    .in_data_7(in_data_7),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N1__width1 muxN_1 (
    .in_data_0(in_data_8),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(3),
    .lo(0),
    .width(4)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(1),
    .lo(0),
    .width(4)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N16__width32 (
    input [31:0] in_data_0,
    input [31:0] in_data_1,
    input [31:0] in_data_10,
    input [31:0] in_data_11,
    input [31:0] in_data_12,
    input [31:0] in_data_13,
    input [31:0] in_data_14,
    input [31:0] in_data_15,
    input [31:0] in_data_2,
    input [31:0] in_data_3,
    input [31:0] in_data_4,
    input [31:0] in_data_5,
    input [31:0] in_data_6,
    input [31:0] in_data_7,
    input [31:0] in_data_8,
    input [31:0] in_data_9,
    input [3:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
wire [31:0] muxN_0_out;
wire [31:0] muxN_1_out;
wire [2:0] sel_slice0_out;
wire [2:0] sel_slice1_out;
coreir_mux #(
    .width(32)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[3]),
    .out(_join_out)
);
commonlib_muxn__N8__width32 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_2(in_data_2),
    .in_data_3(in_data_3),
    .in_data_4(in_data_4),
    .in_data_5(in_data_5),
    .in_data_6(in_data_6),
    .in_data_7(in_data_7),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N8__width32 muxN_1 (
    .in_data_0(in_data_8),
    .in_data_1(in_data_9),
    .in_data_2(in_data_10),
    .in_data_3(in_data_11),
    .in_data_4(in_data_12),
    .in_data_5(in_data_13),
    .in_data_6(in_data_14),
    .in_data_7(in_data_15),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(3),
    .lo(0),
    .width(4)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(3),
    .lo(0),
    .width(4)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N32__width32 (
    input [31:0] in_data_0,
    input [31:0] in_data_1,
    input [31:0] in_data_10,
    input [31:0] in_data_11,
    input [31:0] in_data_12,
    input [31:0] in_data_13,
    input [31:0] in_data_14,
    input [31:0] in_data_15,
    input [31:0] in_data_16,
    input [31:0] in_data_17,
    input [31:0] in_data_18,
    input [31:0] in_data_19,
    input [31:0] in_data_2,
    input [31:0] in_data_20,
    input [31:0] in_data_21,
    input [31:0] in_data_22,
    input [31:0] in_data_23,
    input [31:0] in_data_24,
    input [31:0] in_data_25,
    input [31:0] in_data_26,
    input [31:0] in_data_27,
    input [31:0] in_data_28,
    input [31:0] in_data_29,
    input [31:0] in_data_3,
    input [31:0] in_data_30,
    input [31:0] in_data_31,
    input [31:0] in_data_4,
    input [31:0] in_data_5,
    input [31:0] in_data_6,
    input [31:0] in_data_7,
    input [31:0] in_data_8,
    input [31:0] in_data_9,
    input [4:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
wire [31:0] muxN_0_out;
wire [31:0] muxN_1_out;
wire [3:0] sel_slice0_out;
wire [3:0] sel_slice1_out;
coreir_mux #(
    .width(32)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[4]),
    .out(_join_out)
);
commonlib_muxn__N16__width32 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_10(in_data_10),
    .in_data_11(in_data_11),
    .in_data_12(in_data_12),
    .in_data_13(in_data_13),
    .in_data_14(in_data_14),
    .in_data_15(in_data_15),
    .in_data_2(in_data_2),
    .in_data_3(in_data_3),
    .in_data_4(in_data_4),
    .in_data_5(in_data_5),
    .in_data_6(in_data_6),
    .in_data_7(in_data_7),
    .in_data_8(in_data_8),
    .in_data_9(in_data_9),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N16__width32 muxN_1 (
    .in_data_0(in_data_16),
    .in_data_1(in_data_17),
    .in_data_10(in_data_26),
    .in_data_11(in_data_27),
    .in_data_12(in_data_28),
    .in_data_13(in_data_29),
    .in_data_14(in_data_30),
    .in_data_15(in_data_31),
    .in_data_2(in_data_18),
    .in_data_3(in_data_19),
    .in_data_4(in_data_20),
    .in_data_5(in_data_21),
    .in_data_6(in_data_22),
    .in_data_7(in_data_23),
    .in_data_8(in_data_24),
    .in_data_9(in_data_25),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(4),
    .lo(0),
    .width(5)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(4),
    .lo(0),
    .width(5)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N64__width32 (
    input [31:0] in_data_0,
    input [31:0] in_data_1,
    input [31:0] in_data_10,
    input [31:0] in_data_11,
    input [31:0] in_data_12,
    input [31:0] in_data_13,
    input [31:0] in_data_14,
    input [31:0] in_data_15,
    input [31:0] in_data_16,
    input [31:0] in_data_17,
    input [31:0] in_data_18,
    input [31:0] in_data_19,
    input [31:0] in_data_2,
    input [31:0] in_data_20,
    input [31:0] in_data_21,
    input [31:0] in_data_22,
    input [31:0] in_data_23,
    input [31:0] in_data_24,
    input [31:0] in_data_25,
    input [31:0] in_data_26,
    input [31:0] in_data_27,
    input [31:0] in_data_28,
    input [31:0] in_data_29,
    input [31:0] in_data_3,
    input [31:0] in_data_30,
    input [31:0] in_data_31,
    input [31:0] in_data_32,
    input [31:0] in_data_33,
    input [31:0] in_data_34,
    input [31:0] in_data_35,
    input [31:0] in_data_36,
    input [31:0] in_data_37,
    input [31:0] in_data_38,
    input [31:0] in_data_39,
    input [31:0] in_data_4,
    input [31:0] in_data_40,
    input [31:0] in_data_41,
    input [31:0] in_data_42,
    input [31:0] in_data_43,
    input [31:0] in_data_44,
    input [31:0] in_data_45,
    input [31:0] in_data_46,
    input [31:0] in_data_47,
    input [31:0] in_data_48,
    input [31:0] in_data_49,
    input [31:0] in_data_5,
    input [31:0] in_data_50,
    input [31:0] in_data_51,
    input [31:0] in_data_52,
    input [31:0] in_data_53,
    input [31:0] in_data_54,
    input [31:0] in_data_55,
    input [31:0] in_data_56,
    input [31:0] in_data_57,
    input [31:0] in_data_58,
    input [31:0] in_data_59,
    input [31:0] in_data_6,
    input [31:0] in_data_60,
    input [31:0] in_data_61,
    input [31:0] in_data_62,
    input [31:0] in_data_63,
    input [31:0] in_data_7,
    input [31:0] in_data_8,
    input [31:0] in_data_9,
    input [5:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
wire [31:0] muxN_0_out;
wire [31:0] muxN_1_out;
wire [4:0] sel_slice0_out;
wire [4:0] sel_slice1_out;
coreir_mux #(
    .width(32)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[5]),
    .out(_join_out)
);
commonlib_muxn__N32__width32 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_10(in_data_10),
    .in_data_11(in_data_11),
    .in_data_12(in_data_12),
    .in_data_13(in_data_13),
    .in_data_14(in_data_14),
    .in_data_15(in_data_15),
    .in_data_16(in_data_16),
    .in_data_17(in_data_17),
    .in_data_18(in_data_18),
    .in_data_19(in_data_19),
    .in_data_2(in_data_2),
    .in_data_20(in_data_20),
    .in_data_21(in_data_21),
    .in_data_22(in_data_22),
    .in_data_23(in_data_23),
    .in_data_24(in_data_24),
    .in_data_25(in_data_25),
    .in_data_26(in_data_26),
    .in_data_27(in_data_27),
    .in_data_28(in_data_28),
    .in_data_29(in_data_29),
    .in_data_3(in_data_3),
    .in_data_30(in_data_30),
    .in_data_31(in_data_31),
    .in_data_4(in_data_4),
    .in_data_5(in_data_5),
    .in_data_6(in_data_6),
    .in_data_7(in_data_7),
    .in_data_8(in_data_8),
    .in_data_9(in_data_9),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N32__width32 muxN_1 (
    .in_data_0(in_data_32),
    .in_data_1(in_data_33),
    .in_data_10(in_data_42),
    .in_data_11(in_data_43),
    .in_data_12(in_data_44),
    .in_data_13(in_data_45),
    .in_data_14(in_data_46),
    .in_data_15(in_data_47),
    .in_data_16(in_data_48),
    .in_data_17(in_data_49),
    .in_data_18(in_data_50),
    .in_data_19(in_data_51),
    .in_data_2(in_data_34),
    .in_data_20(in_data_52),
    .in_data_21(in_data_53),
    .in_data_22(in_data_54),
    .in_data_23(in_data_55),
    .in_data_24(in_data_56),
    .in_data_25(in_data_57),
    .in_data_26(in_data_58),
    .in_data_27(in_data_59),
    .in_data_28(in_data_60),
    .in_data_29(in_data_61),
    .in_data_3(in_data_35),
    .in_data_30(in_data_62),
    .in_data_31(in_data_63),
    .in_data_4(in_data_36),
    .in_data_5(in_data_37),
    .in_data_6(in_data_38),
    .in_data_7(in_data_39),
    .in_data_8(in_data_40),
    .in_data_9(in_data_41),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(5),
    .lo(0),
    .width(6)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(5),
    .lo(0),
    .width(6)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N20__width32 (
    input [31:0] in_data_0,
    input [31:0] in_data_1,
    input [31:0] in_data_10,
    input [31:0] in_data_11,
    input [31:0] in_data_12,
    input [31:0] in_data_13,
    input [31:0] in_data_14,
    input [31:0] in_data_15,
    input [31:0] in_data_16,
    input [31:0] in_data_17,
    input [31:0] in_data_18,
    input [31:0] in_data_19,
    input [31:0] in_data_2,
    input [31:0] in_data_3,
    input [31:0] in_data_4,
    input [31:0] in_data_5,
    input [31:0] in_data_6,
    input [31:0] in_data_7,
    input [31:0] in_data_8,
    input [31:0] in_data_9,
    input [4:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
wire [31:0] muxN_0_out;
wire [31:0] muxN_1_out;
wire [3:0] sel_slice0_out;
wire [1:0] sel_slice1_out;
coreir_mux #(
    .width(32)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[4]),
    .out(_join_out)
);
commonlib_muxn__N16__width32 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_10(in_data_10),
    .in_data_11(in_data_11),
    .in_data_12(in_data_12),
    .in_data_13(in_data_13),
    .in_data_14(in_data_14),
    .in_data_15(in_data_15),
    .in_data_2(in_data_2),
    .in_data_3(in_data_3),
    .in_data_4(in_data_4),
    .in_data_5(in_data_5),
    .in_data_6(in_data_6),
    .in_data_7(in_data_7),
    .in_data_8(in_data_8),
    .in_data_9(in_data_9),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N4__width32 muxN_1 (
    .in_data_0(in_data_16),
    .in_data_1(in_data_17),
    .in_data_2(in_data_18),
    .in_data_3(in_data_19),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(4),
    .lo(0),
    .width(5)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(2),
    .lo(0),
    .width(5)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N84__width32 (
    input [31:0] in_data_0,
    input [31:0] in_data_1,
    input [31:0] in_data_10,
    input [31:0] in_data_11,
    input [31:0] in_data_12,
    input [31:0] in_data_13,
    input [31:0] in_data_14,
    input [31:0] in_data_15,
    input [31:0] in_data_16,
    input [31:0] in_data_17,
    input [31:0] in_data_18,
    input [31:0] in_data_19,
    input [31:0] in_data_2,
    input [31:0] in_data_20,
    input [31:0] in_data_21,
    input [31:0] in_data_22,
    input [31:0] in_data_23,
    input [31:0] in_data_24,
    input [31:0] in_data_25,
    input [31:0] in_data_26,
    input [31:0] in_data_27,
    input [31:0] in_data_28,
    input [31:0] in_data_29,
    input [31:0] in_data_3,
    input [31:0] in_data_30,
    input [31:0] in_data_31,
    input [31:0] in_data_32,
    input [31:0] in_data_33,
    input [31:0] in_data_34,
    input [31:0] in_data_35,
    input [31:0] in_data_36,
    input [31:0] in_data_37,
    input [31:0] in_data_38,
    input [31:0] in_data_39,
    input [31:0] in_data_4,
    input [31:0] in_data_40,
    input [31:0] in_data_41,
    input [31:0] in_data_42,
    input [31:0] in_data_43,
    input [31:0] in_data_44,
    input [31:0] in_data_45,
    input [31:0] in_data_46,
    input [31:0] in_data_47,
    input [31:0] in_data_48,
    input [31:0] in_data_49,
    input [31:0] in_data_5,
    input [31:0] in_data_50,
    input [31:0] in_data_51,
    input [31:0] in_data_52,
    input [31:0] in_data_53,
    input [31:0] in_data_54,
    input [31:0] in_data_55,
    input [31:0] in_data_56,
    input [31:0] in_data_57,
    input [31:0] in_data_58,
    input [31:0] in_data_59,
    input [31:0] in_data_6,
    input [31:0] in_data_60,
    input [31:0] in_data_61,
    input [31:0] in_data_62,
    input [31:0] in_data_63,
    input [31:0] in_data_64,
    input [31:0] in_data_65,
    input [31:0] in_data_66,
    input [31:0] in_data_67,
    input [31:0] in_data_68,
    input [31:0] in_data_69,
    input [31:0] in_data_7,
    input [31:0] in_data_70,
    input [31:0] in_data_71,
    input [31:0] in_data_72,
    input [31:0] in_data_73,
    input [31:0] in_data_74,
    input [31:0] in_data_75,
    input [31:0] in_data_76,
    input [31:0] in_data_77,
    input [31:0] in_data_78,
    input [31:0] in_data_79,
    input [31:0] in_data_8,
    input [31:0] in_data_80,
    input [31:0] in_data_81,
    input [31:0] in_data_82,
    input [31:0] in_data_83,
    input [31:0] in_data_9,
    input [6:0] in_sel,
    output [31:0] out
);
wire [31:0] _join_out;
wire [31:0] muxN_0_out;
wire [31:0] muxN_1_out;
wire [5:0] sel_slice0_out;
wire [4:0] sel_slice1_out;
coreir_mux #(
    .width(32)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[6]),
    .out(_join_out)
);
commonlib_muxn__N64__width32 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_10(in_data_10),
    .in_data_11(in_data_11),
    .in_data_12(in_data_12),
    .in_data_13(in_data_13),
    .in_data_14(in_data_14),
    .in_data_15(in_data_15),
    .in_data_16(in_data_16),
    .in_data_17(in_data_17),
    .in_data_18(in_data_18),
    .in_data_19(in_data_19),
    .in_data_2(in_data_2),
    .in_data_20(in_data_20),
    .in_data_21(in_data_21),
    .in_data_22(in_data_22),
    .in_data_23(in_data_23),
    .in_data_24(in_data_24),
    .in_data_25(in_data_25),
    .in_data_26(in_data_26),
    .in_data_27(in_data_27),
    .in_data_28(in_data_28),
    .in_data_29(in_data_29),
    .in_data_3(in_data_3),
    .in_data_30(in_data_30),
    .in_data_31(in_data_31),
    .in_data_32(in_data_32),
    .in_data_33(in_data_33),
    .in_data_34(in_data_34),
    .in_data_35(in_data_35),
    .in_data_36(in_data_36),
    .in_data_37(in_data_37),
    .in_data_38(in_data_38),
    .in_data_39(in_data_39),
    .in_data_4(in_data_4),
    .in_data_40(in_data_40),
    .in_data_41(in_data_41),
    .in_data_42(in_data_42),
    .in_data_43(in_data_43),
    .in_data_44(in_data_44),
    .in_data_45(in_data_45),
    .in_data_46(in_data_46),
    .in_data_47(in_data_47),
    .in_data_48(in_data_48),
    .in_data_49(in_data_49),
    .in_data_5(in_data_5),
    .in_data_50(in_data_50),
    .in_data_51(in_data_51),
    .in_data_52(in_data_52),
    .in_data_53(in_data_53),
    .in_data_54(in_data_54),
    .in_data_55(in_data_55),
    .in_data_56(in_data_56),
    .in_data_57(in_data_57),
    .in_data_58(in_data_58),
    .in_data_59(in_data_59),
    .in_data_6(in_data_6),
    .in_data_60(in_data_60),
    .in_data_61(in_data_61),
    .in_data_62(in_data_62),
    .in_data_63(in_data_63),
    .in_data_7(in_data_7),
    .in_data_8(in_data_8),
    .in_data_9(in_data_9),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N20__width32 muxN_1 (
    .in_data_0(in_data_64),
    .in_data_1(in_data_65),
    .in_data_10(in_data_74),
    .in_data_11(in_data_75),
    .in_data_12(in_data_76),
    .in_data_13(in_data_77),
    .in_data_14(in_data_78),
    .in_data_15(in_data_79),
    .in_data_16(in_data_80),
    .in_data_17(in_data_81),
    .in_data_18(in_data_82),
    .in_data_19(in_data_83),
    .in_data_2(in_data_66),
    .in_data_3(in_data_67),
    .in_data_4(in_data_68),
    .in_data_5(in_data_69),
    .in_data_6(in_data_70),
    .in_data_7(in_data_71),
    .in_data_8(in_data_72),
    .in_data_9(in_data_73),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(6),
    .lo(0),
    .width(7)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(5),
    .lo(0),
    .width(7)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N16__width16 (
    input [15:0] in_data_0,
    input [15:0] in_data_1,
    input [15:0] in_data_10,
    input [15:0] in_data_11,
    input [15:0] in_data_12,
    input [15:0] in_data_13,
    input [15:0] in_data_14,
    input [15:0] in_data_15,
    input [15:0] in_data_2,
    input [15:0] in_data_3,
    input [15:0] in_data_4,
    input [15:0] in_data_5,
    input [15:0] in_data_6,
    input [15:0] in_data_7,
    input [15:0] in_data_8,
    input [15:0] in_data_9,
    input [3:0] in_sel,
    output [15:0] out
);
wire [15:0] _join_out;
wire [15:0] muxN_0_out;
wire [15:0] muxN_1_out;
wire [2:0] sel_slice0_out;
wire [2:0] sel_slice1_out;
coreir_mux #(
    .width(16)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[3]),
    .out(_join_out)
);
commonlib_muxn__N8__width16 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_2(in_data_2),
    .in_data_3(in_data_3),
    .in_data_4(in_data_4),
    .in_data_5(in_data_5),
    .in_data_6(in_data_6),
    .in_data_7(in_data_7),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N8__width16 muxN_1 (
    .in_data_0(in_data_8),
    .in_data_1(in_data_9),
    .in_data_2(in_data_10),
    .in_data_3(in_data_11),
    .in_data_4(in_data_12),
    .in_data_5(in_data_13),
    .in_data_6(in_data_14),
    .in_data_7(in_data_15),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(3),
    .lo(0),
    .width(4)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(3),
    .lo(0),
    .width(4)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N20__width16 (
    input [15:0] in_data_0,
    input [15:0] in_data_1,
    input [15:0] in_data_10,
    input [15:0] in_data_11,
    input [15:0] in_data_12,
    input [15:0] in_data_13,
    input [15:0] in_data_14,
    input [15:0] in_data_15,
    input [15:0] in_data_16,
    input [15:0] in_data_17,
    input [15:0] in_data_18,
    input [15:0] in_data_19,
    input [15:0] in_data_2,
    input [15:0] in_data_3,
    input [15:0] in_data_4,
    input [15:0] in_data_5,
    input [15:0] in_data_6,
    input [15:0] in_data_7,
    input [15:0] in_data_8,
    input [15:0] in_data_9,
    input [4:0] in_sel,
    output [15:0] out
);
wire [15:0] _join_out;
wire [15:0] muxN_0_out;
wire [15:0] muxN_1_out;
wire [3:0] sel_slice0_out;
wire [1:0] sel_slice1_out;
coreir_mux #(
    .width(16)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[4]),
    .out(_join_out)
);
commonlib_muxn__N16__width16 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_10(in_data_10),
    .in_data_11(in_data_11),
    .in_data_12(in_data_12),
    .in_data_13(in_data_13),
    .in_data_14(in_data_14),
    .in_data_15(in_data_15),
    .in_data_2(in_data_2),
    .in_data_3(in_data_3),
    .in_data_4(in_data_4),
    .in_data_5(in_data_5),
    .in_data_6(in_data_6),
    .in_data_7(in_data_7),
    .in_data_8(in_data_8),
    .in_data_9(in_data_9),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N4__width16 muxN_1 (
    .in_data_0(in_data_16),
    .in_data_1(in_data_17),
    .in_data_2(in_data_18),
    .in_data_3(in_data_19),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(4),
    .lo(0),
    .width(5)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(2),
    .lo(0),
    .width(5)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N16__width1 (
    input [0:0] in_data_0,
    input [0:0] in_data_1,
    input [0:0] in_data_10,
    input [0:0] in_data_11,
    input [0:0] in_data_12,
    input [0:0] in_data_13,
    input [0:0] in_data_14,
    input [0:0] in_data_15,
    input [0:0] in_data_2,
    input [0:0] in_data_3,
    input [0:0] in_data_4,
    input [0:0] in_data_5,
    input [0:0] in_data_6,
    input [0:0] in_data_7,
    input [0:0] in_data_8,
    input [0:0] in_data_9,
    input [3:0] in_sel,
    output [0:0] out
);
wire [0:0] _join_out;
wire [0:0] muxN_0_out;
wire [0:0] muxN_1_out;
wire [2:0] sel_slice0_out;
wire [2:0] sel_slice1_out;
coreir_mux #(
    .width(1)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[3]),
    .out(_join_out)
);
commonlib_muxn__N8__width1 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_2(in_data_2),
    .in_data_3(in_data_3),
    .in_data_4(in_data_4),
    .in_data_5(in_data_5),
    .in_data_6(in_data_6),
    .in_data_7(in_data_7),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N8__width1 muxN_1 (
    .in_data_0(in_data_8),
    .in_data_1(in_data_9),
    .in_data_2(in_data_10),
    .in_data_3(in_data_11),
    .in_data_4(in_data_12),
    .in_data_5(in_data_13),
    .in_data_6(in_data_14),
    .in_data_7(in_data_15),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(3),
    .lo(0),
    .width(4)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(3),
    .lo(0),
    .width(4)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module commonlib_muxn__N20__width1 (
    input [0:0] in_data_0,
    input [0:0] in_data_1,
    input [0:0] in_data_10,
    input [0:0] in_data_11,
    input [0:0] in_data_12,
    input [0:0] in_data_13,
    input [0:0] in_data_14,
    input [0:0] in_data_15,
    input [0:0] in_data_16,
    input [0:0] in_data_17,
    input [0:0] in_data_18,
    input [0:0] in_data_19,
    input [0:0] in_data_2,
    input [0:0] in_data_3,
    input [0:0] in_data_4,
    input [0:0] in_data_5,
    input [0:0] in_data_6,
    input [0:0] in_data_7,
    input [0:0] in_data_8,
    input [0:0] in_data_9,
    input [4:0] in_sel,
    output [0:0] out
);
wire [0:0] _join_out;
wire [0:0] muxN_0_out;
wire [0:0] muxN_1_out;
wire [3:0] sel_slice0_out;
wire [1:0] sel_slice1_out;
coreir_mux #(
    .width(1)
) _join (
    .in0(muxN_0_out),
    .in1(muxN_1_out),
    .sel(in_sel[4]),
    .out(_join_out)
);
commonlib_muxn__N16__width1 muxN_0 (
    .in_data_0(in_data_0),
    .in_data_1(in_data_1),
    .in_data_10(in_data_10),
    .in_data_11(in_data_11),
    .in_data_12(in_data_12),
    .in_data_13(in_data_13),
    .in_data_14(in_data_14),
    .in_data_15(in_data_15),
    .in_data_2(in_data_2),
    .in_data_3(in_data_3),
    .in_data_4(in_data_4),
    .in_data_5(in_data_5),
    .in_data_6(in_data_6),
    .in_data_7(in_data_7),
    .in_data_8(in_data_8),
    .in_data_9(in_data_9),
    .in_sel(sel_slice0_out),
    .out(muxN_0_out)
);
commonlib_muxn__N4__width1 muxN_1 (
    .in_data_0(in_data_16),
    .in_data_1(in_data_17),
    .in_data_2(in_data_18),
    .in_data_3(in_data_19),
    .in_sel(sel_slice1_out),
    .out(muxN_1_out)
);
coreir_slice #(
    .hi(4),
    .lo(0),
    .width(5)
) sel_slice0 (
    .in(in_sel),
    .out(sel_slice0_out)
);
coreir_slice #(
    .hi(2),
    .lo(0),
    .width(5)
) sel_slice1 (
    .in(in_sel),
    .out(sel_slice1_out)
);
assign out = _join_out;
endmodule

module chain_chain_en (
    input [22:0] I,
    output [0:0] O
);
assign O = I[0];
endmodule

module SUB (
    input [15:0] a,
    input [15:0] b,
    output [15:0] O0,
    output O1,
    output O2,
    output O3,
    output O4,
    output O5,
    input CLK,
    input ASYNCRESET
);
wire bit_const_0_None_out;
wire [15:0] const_0_16_out;
wire [16:0] const_1_17_out;
wire magma_Bit_and_inst0_out;
wire magma_Bit_and_inst1_out;
wire magma_Bit_and_inst2_out;
wire magma_Bit_and_inst3_out;
wire magma_Bit_not_inst0_out;
wire magma_Bit_not_inst1_out;
wire magma_Bit_not_inst2_out;
wire magma_Bit_or_inst0_out;
wire magma_Bits_16_eq_inst0_out;
wire [15:0] magma_Bits_16_not_inst0_out;
wire [16:0] magma_Bits_17_add_inst0_out;
wire [16:0] magma_Bits_17_add_inst1_out;
corebit_const #(
    .value(1'b0)
) bit_const_0_None (
    .out(bit_const_0_None_out)
);
coreir_const #(
    .value(16'h0000),
    .width(16)
) const_0_16 (
    .out(const_0_16_out)
);
coreir_const #(
    .value(17'h00001),
    .width(17)
) const_1_17 (
    .out(const_1_17_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(a[15]),
    .in1(magma_Bits_16_not_inst0_out[15]),
    .out(magma_Bit_and_inst0_out)
);
corebit_and magma_Bit_and_inst1 (
    .in0(magma_Bit_and_inst0_out),
    .in1(magma_Bit_not_inst0_out),
    .out(magma_Bit_and_inst1_out)
);
corebit_and magma_Bit_and_inst2 (
    .in0(magma_Bit_not_inst1_out),
    .in1(magma_Bit_not_inst2_out),
    .out(magma_Bit_and_inst2_out)
);
corebit_and magma_Bit_and_inst3 (
    .in0(magma_Bit_and_inst2_out),
    .in1(magma_Bits_17_add_inst1_out[15]),
    .out(magma_Bit_and_inst3_out)
);
corebit_not magma_Bit_not_inst0 (
    .in(magma_Bits_17_add_inst1_out[15]),
    .out(magma_Bit_not_inst0_out)
);
corebit_not magma_Bit_not_inst1 (
    .in(a[15]),
    .out(magma_Bit_not_inst1_out)
);
corebit_not magma_Bit_not_inst2 (
    .in(magma_Bits_16_not_inst0_out[15]),
    .out(magma_Bit_not_inst2_out)
);
corebit_or magma_Bit_or_inst0 (
    .in0(magma_Bit_and_inst1_out),
    .in1(magma_Bit_and_inst3_out),
    .out(magma_Bit_or_inst0_out)
);
coreir_eq #(
    .width(16)
) magma_Bits_16_eq_inst0 (
    .in0(magma_Bits_17_add_inst1_out[15:0]),
    .in1(const_0_16_out),
    .out(magma_Bits_16_eq_inst0_out)
);
coreir_not #(
    .width(16)
) magma_Bits_16_not_inst0 (
    .in(b),
    .out(magma_Bits_16_not_inst0_out)
);
wire [16:0] magma_Bits_17_add_inst0_in0;
assign magma_Bits_17_add_inst0_in0 = {bit_const_0_None_out,a[15:0]};
wire [16:0] magma_Bits_17_add_inst0_in1;
assign magma_Bits_17_add_inst0_in1 = {bit_const_0_None_out,magma_Bits_16_not_inst0_out[15:0]};
coreir_add #(
    .width(17)
) magma_Bits_17_add_inst0 (
    .in0(magma_Bits_17_add_inst0_in0),
    .in1(magma_Bits_17_add_inst0_in1),
    .out(magma_Bits_17_add_inst0_out)
);
coreir_add #(
    .width(17)
) magma_Bits_17_add_inst1 (
    .in0(magma_Bits_17_add_inst0_out),
    .in1(const_1_17_out),
    .out(magma_Bits_17_add_inst1_out)
);
assign O0 = magma_Bits_17_add_inst1_out[15:0];
assign O1 = magma_Bits_17_add_inst1_out[16];
assign O2 = magma_Bits_16_eq_inst0_out;
assign O3 = magma_Bits_17_add_inst1_out[15];
assign O4 = magma_Bits_17_add_inst1_out[16];
assign O5 = magma_Bit_or_inst0_out;
endmodule

module SHR (
    input [0:0] signed_,
    input [15:0] a,
    input [15:0] b,
    output [15:0] O0,
    output O1,
    output O2,
    output O3,
    output O4,
    output O5,
    input CLK,
    input ASYNCRESET
);
wire [15:0] Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire bit_const_0_None_out;
wire [15:0] const_0_16_out;
wire [0:0] const_1_1_out;
wire [15:0] magma_Bits_16_ashr_inst0_out;
wire magma_Bits_16_eq_inst0_out;
wire [15:0] magma_Bits_16_lshr_inst0_out;
wire magma_Bits_1_eq_inst0_out;
coreir_mux #(
    .width(16)
) Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(magma_Bits_16_lshr_inst0_out),
    .in1(magma_Bits_16_ashr_inst0_out),
    .sel(magma_Bits_1_eq_inst0_out),
    .out(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
corebit_const #(
    .value(1'b0)
) bit_const_0_None (
    .out(bit_const_0_None_out)
);
coreir_const #(
    .value(16'h0000),
    .width(16)
) const_0_16 (
    .out(const_0_16_out)
);
coreir_const #(
    .value(1'h1),
    .width(1)
) const_1_1 (
    .out(const_1_1_out)
);
coreir_ashr #(
    .width(16)
) magma_Bits_16_ashr_inst0 (
    .in0(a),
    .in1(b),
    .out(magma_Bits_16_ashr_inst0_out)
);
coreir_eq #(
    .width(16)
) magma_Bits_16_eq_inst0 (
    .in0(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(const_0_16_out),
    .out(magma_Bits_16_eq_inst0_out)
);
coreir_lshr #(
    .width(16)
) magma_Bits_16_lshr_inst0 (
    .in0(a),
    .in1(b),
    .out(magma_Bits_16_lshr_inst0_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst0 (
    .in0(signed_),
    .in1(const_1_1_out),
    .out(magma_Bits_1_eq_inst0_out)
);
assign O0 = Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign O1 = bit_const_0_None_out;
assign O2 = magma_Bits_16_eq_inst0_out;
assign O3 = Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out[15];
assign O4 = bit_const_0_None_out;
assign O5 = bit_const_0_None_out;
endmodule

module SB_T4_WEST_SB_OUT_B1_sel_unq1 (
    input [3:0] I,
    output [3:0] O
);
assign O = I;
endmodule

module SB_T4_WEST_SB_OUT_B1_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[27:26];
endmodule

module SB_T4_WEST_SB_OUT_B16_sel_unq1 (
    input [17:0] I,
    output [2:0] O
);
assign O = I[17:15];
endmodule

module SB_T4_WEST_SB_OUT_B16_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[27:26];
endmodule

module SB_T4_SOUTH_SB_OUT_B1_sel_unq1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[31:28];
endmodule

module SB_T4_SOUTH_SB_OUT_B1_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[25:24];
endmodule

module SB_T4_SOUTH_SB_OUT_B16_sel_unq1 (
    input [17:0] I,
    output [2:0] O
);
assign O = I[14:12];
endmodule

module SB_T4_SOUTH_SB_OUT_B16_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[25:24];
endmodule

module SB_T4_NORTH_SB_OUT_B1_sel_unq1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[27:24];
endmodule

module SB_T4_NORTH_SB_OUT_B1_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[23:22];
endmodule

module SB_T4_NORTH_SB_OUT_B16_sel_unq1 (
    input [17:0] I,
    output [2:0] O
);
assign O = I[11:9];
endmodule

module SB_T4_NORTH_SB_OUT_B16_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[23:22];
endmodule

module SB_T4_EAST_SB_OUT_B1_sel_unq1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[23:20];
endmodule

module SB_T4_EAST_SB_OUT_B1_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[21:20];
endmodule

module SB_T4_EAST_SB_OUT_B16_sel_unq1 (
    input [17:0] I,
    output [2:0] O
);
assign O = I[8:6];
endmodule

module SB_T4_EAST_SB_OUT_B16_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[21:20];
endmodule

module SB_T3_WEST_SB_OUT_B1_sel_unq1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[19:16];
endmodule

module SB_T3_WEST_SB_OUT_B1_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[19:18];
endmodule

module SB_T3_WEST_SB_OUT_B16_sel_unq1 (
    input [17:0] I,
    output [2:0] O
);
assign O = I[5:3];
endmodule

module SB_T3_WEST_SB_OUT_B16_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[19:18];
endmodule

module SB_T3_SOUTH_SB_OUT_B1_sel_unq1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[15:12];
endmodule

module SB_T3_SOUTH_SB_OUT_B1_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[17:16];
endmodule

module SB_T3_SOUTH_SB_OUT_B16_sel_unq1 (
    input [17:0] I,
    output [2:0] O
);
assign O = I[2:0];
endmodule

module SB_T3_SOUTH_SB_OUT_B16_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[17:16];
endmodule

module SB_T3_NORTH_SB_OUT_B1_sel_unq1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[11:8];
endmodule

module SB_T3_NORTH_SB_OUT_B1_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[15:14];
endmodule

module SB_T3_NORTH_SB_OUT_B16_sel_unq1 (
    input [29:0] I,
    output [2:0] O
);
assign O = I[29:27];
endmodule

module SB_T3_NORTH_SB_OUT_B16_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[15:14];
endmodule

module SB_T3_EAST_SB_OUT_B1_sel_unq1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[7:4];
endmodule

module SB_T3_EAST_SB_OUT_B1_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[13:12];
endmodule

module SB_T3_EAST_SB_OUT_B16_sel_unq1 (
    input [29:0] I,
    output [2:0] O
);
assign O = I[26:24];
endmodule

module SB_T3_EAST_SB_OUT_B16_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[13:12];
endmodule

module SB_T2_WEST_SB_OUT_B1_sel_unq1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module SB_T2_WEST_SB_OUT_B1_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[11:10];
endmodule

module SB_T2_WEST_SB_OUT_B16_sel_unq1 (
    input [29:0] I,
    output [2:0] O
);
assign O = I[23:21];
endmodule

module SB_T2_WEST_SB_OUT_B16_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[11:10];
endmodule

module SB_T2_SOUTH_SB_OUT_B1_sel_unq1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[31:28];
endmodule

module SB_T2_SOUTH_SB_OUT_B1_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[9:8];
endmodule

module SB_T2_SOUTH_SB_OUT_B16_sel_unq1 (
    input [29:0] I,
    output [2:0] O
);
assign O = I[20:18];
endmodule

module SB_T2_SOUTH_SB_OUT_B16_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[9:8];
endmodule

module SB_T2_NORTH_SB_OUT_B1_sel_unq1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[27:24];
endmodule

module SB_T2_NORTH_SB_OUT_B1_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[7:6];
endmodule

module SB_T2_NORTH_SB_OUT_B16_sel_unq1 (
    input [29:0] I,
    output [2:0] O
);
assign O = I[17:15];
endmodule

module SB_T2_NORTH_SB_OUT_B16_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[7:6];
endmodule

module SB_T2_EAST_SB_OUT_B1_sel_unq1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[23:20];
endmodule

module SB_T2_EAST_SB_OUT_B1_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[5:4];
endmodule

module SB_T2_EAST_SB_OUT_B16_sel_unq1 (
    input [29:0] I,
    output [2:0] O
);
assign O = I[14:12];
endmodule

module SB_T2_EAST_SB_OUT_B16_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[5:4];
endmodule

module SB_T1_WEST_SB_OUT_B1_sel_unq1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[19:16];
endmodule

module SB_T1_WEST_SB_OUT_B1_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[3:2];
endmodule

module SB_T1_WEST_SB_OUT_B16_sel_unq1 (
    input [29:0] I,
    output [2:0] O
);
assign O = I[11:9];
endmodule

module SB_T1_WEST_SB_OUT_B16_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[3:2];
endmodule

module SB_T1_SOUTH_SB_OUT_B1_sel_unq1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[15:12];
endmodule

module SB_T1_SOUTH_SB_OUT_B1_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[1:0];
endmodule

module SB_T1_SOUTH_SB_OUT_B16_sel_unq1 (
    input [29:0] I,
    output [2:0] O
);
assign O = I[8:6];
endmodule

module SB_T1_SOUTH_SB_OUT_B16_sel (
    input [27:0] I,
    output [1:0] O
);
assign O = I[1:0];
endmodule

module SB_T1_NORTH_SB_OUT_B1_sel_unq1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[11:8];
endmodule

module SB_T1_NORTH_SB_OUT_B1_sel (
    input [31:0] I,
    output [1:0] O
);
assign O = I[31:30];
endmodule

module SB_T1_NORTH_SB_OUT_B16_sel_unq1 (
    input [29:0] I,
    output [2:0] O
);
assign O = I[5:3];
endmodule

module SB_T1_NORTH_SB_OUT_B16_sel (
    input [31:0] I,
    output [1:0] O
);
assign O = I[31:30];
endmodule

module SB_T1_EAST_SB_OUT_B1_sel_unq1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[7:4];
endmodule

module SB_T1_EAST_SB_OUT_B1_sel (
    input [31:0] I,
    output [1:0] O
);
assign O = I[29:28];
endmodule

module SB_T1_EAST_SB_OUT_B16_sel_unq1 (
    input [29:0] I,
    output [2:0] O
);
assign O = I[2:0];
endmodule

module SB_T1_EAST_SB_OUT_B16_sel (
    input [31:0] I,
    output [1:0] O
);
assign O = I[29:28];
endmodule

module SB_T0_WEST_SB_OUT_B1_sel_unq1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[3:0];
endmodule

module SB_T0_WEST_SB_OUT_B1_sel (
    input [31:0] I,
    output [1:0] O
);
assign O = I[27:26];
endmodule

module SB_T0_WEST_SB_OUT_B16_sel_unq1 (
    input [31:0] I,
    output [2:0] O
);
assign O = I[31:29];
endmodule

module SB_T0_WEST_SB_OUT_B16_sel (
    input [31:0] I,
    output [1:0] O
);
assign O = I[27:26];
endmodule

module SB_T0_SOUTH_SB_OUT_B1_sel_unq1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[31:28];
endmodule

module SB_T0_SOUTH_SB_OUT_B1_sel (
    input [31:0] I,
    output [1:0] O
);
assign O = I[25:24];
endmodule

module SB_T0_SOUTH_SB_OUT_B16_sel_unq1 (
    input [31:0] I,
    output [2:0] O
);
assign O = I[28:26];
endmodule

module SB_T0_SOUTH_SB_OUT_B16_sel (
    input [31:0] I,
    output [1:0] O
);
assign O = I[25:24];
endmodule

module SB_T0_NORTH_SB_OUT_B1_sel_unq1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[27:24];
endmodule

module SB_T0_NORTH_SB_OUT_B1_sel (
    input [31:0] I,
    output [1:0] O
);
assign O = I[23:22];
endmodule

module SB_T0_NORTH_SB_OUT_B16_sel_unq1 (
    input [31:0] I,
    output [2:0] O
);
assign O = I[25:23];
endmodule

module SB_T0_NORTH_SB_OUT_B16_sel (
    input [31:0] I,
    output [1:0] O
);
assign O = I[23:22];
endmodule

module SB_T0_EAST_SB_OUT_B1_sel_unq1 (
    input [31:0] I,
    output [3:0] O
);
assign O = I[23:20];
endmodule

module SB_T0_EAST_SB_OUT_B1_sel (
    input [31:0] I,
    output [1:0] O
);
assign O = I[21:20];
endmodule

module SB_T0_EAST_SB_OUT_B16_sel_unq1 (
    input [31:0] I,
    output [2:0] O
);
assign O = I[22:20];
endmodule

module SB_T0_EAST_SB_OUT_B16_sel (
    input [31:0] I,
    output [1:0] O
);
assign O = I[21:20];
endmodule

module Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_5 (
    input [4:0] I,
    output [4:0] O,
    input CLK,
    input CE,
    input ASYNCRESET
);
wire [4:0] value__CE_out;
regCE_arst #(
    .init(5'h00),
    .width(5)
) value__CE (
    .in(I),
    .ce(CE),
    .out(value__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = value__CE_out;
endmodule

module Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_4 (
    input [3:0] I,
    output [3:0] O,
    input CLK,
    input CE,
    input ASYNCRESET
);
wire [3:0] value__CE_out;
regCE_arst #(
    .init(4'h0),
    .width(4)
) value__CE (
    .in(I),
    .ce(CE),
    .out(value__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = value__CE_out;
endmodule

module Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 (
    input [31:0] I,
    output [31:0] O,
    input CLK,
    input CE,
    input ASYNCRESET
);
wire [31:0] value__CE_out;
regCE_arst #(
    .init(32'h00000000),
    .width(32)
) value__CE (
    .in(I),
    .ce(CE),
    .out(value__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = value__CE_out;
endmodule

module Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_31 (
    input [30:0] I,
    output [30:0] O,
    input CLK,
    input CE,
    input ASYNCRESET
);
wire [30:0] value__CE_out;
regCE_arst #(
    .init(31'h00000000),
    .width(31)
) value__CE (
    .in(I),
    .ce(CE),
    .out(value__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = value__CE_out;
endmodule

module Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_30 (
    input [29:0] I,
    output [29:0] O,
    input CLK,
    input CE,
    input ASYNCRESET
);
wire [29:0] value__CE_out;
regCE_arst #(
    .init(30'h00000000),
    .width(30)
) value__CE (
    .in(I),
    .ce(CE),
    .out(value__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = value__CE_out;
endmodule

module Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_29 (
    input [28:0] I,
    output [28:0] O,
    input CLK,
    input CE,
    input ASYNCRESET
);
wire [28:0] value__CE_out;
regCE_arst #(
    .init(29'h00000000),
    .width(29)
) value__CE (
    .in(I),
    .ce(CE),
    .out(value__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = value__CE_out;
endmodule

module Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_28 (
    input [27:0] I,
    output [27:0] O,
    input CLK,
    input CE,
    input ASYNCRESET
);
wire [27:0] value__CE_out;
regCE_arst #(
    .init(28'h0000000),
    .width(28)
) value__CE (
    .in(I),
    .ce(CE),
    .out(value__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = value__CE_out;
endmodule

module Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27 (
    input [26:0] I,
    output [26:0] O,
    input CLK,
    input CE,
    input ASYNCRESET
);
wire [26:0] value__CE_out;
regCE_arst #(
    .init(27'h0000000),
    .width(27)
) value__CE (
    .in(I),
    .ce(CE),
    .out(value__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = value__CE_out;
endmodule

module Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_25 (
    input [24:0] I,
    output [24:0] O,
    input CLK,
    input CE,
    input ASYNCRESET
);
wire [24:0] value__CE_out;
regCE_arst #(
    .init(25'h0000000),
    .width(25)
) value__CE (
    .in(I),
    .ce(CE),
    .out(value__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = value__CE_out;
endmodule

module Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_23 (
    input [22:0] I,
    output [22:0] O,
    input CLK,
    input CE,
    input ASYNCRESET
);
wire [22:0] value__CE_out;
regCE_arst #(
    .init(23'h000000),
    .width(23)
) value__CE (
    .in(I),
    .ce(CE),
    .out(value__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = value__CE_out;
endmodule

module Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20 (
    input [19:0] I,
    output [19:0] O,
    input CLK,
    input CE,
    input ASYNCRESET
);
wire [19:0] value__CE_out;
regCE_arst #(
    .init(20'h00000),
    .width(20)
) value__CE (
    .in(I),
    .ce(CE),
    .out(value__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = value__CE_out;
endmodule

module Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_18 (
    input [17:0] I,
    output [17:0] O,
    input CLK,
    input CE,
    input ASYNCRESET
);
wire [17:0] value__CE_out;
regCE_arst #(
    .init(18'h00000),
    .width(18)
) value__CE (
    .in(I),
    .ce(CE),
    .out(value__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = value__CE_out;
endmodule

module Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17 (
    input [16:0] I,
    output [16:0] O,
    input CLK,
    input CE,
    input ASYNCRESET
);
wire [16:0] value__CE_out;
regCE_arst #(
    .init(17'h00000),
    .width(17)
) value__CE (
    .in(I),
    .ce(CE),
    .out(value__CE_out),
    .clk(CLK),
    .arst(ASYNCRESET)
);
assign O = value__CE_out;
endmodule

module Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 (
    input [15:0] I,
    output [15:0] O,
    input CLK,
    input CE
);
wire [15:0] value__CE_out;
regCE #(
    .width(16)
) value__CE (
    .in(I),
    .ce(CE),
    .out(value__CE_out),
    .clk(CLK)
);
assign O = value__CE_out;
endmodule

module Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 (
    input [0:0] I,
    output [0:0] O,
    input CLK,
    input CE
);
wire [0:0] value__CE_out;
regCE #(
    .width(1)
) value__CE (
    .in(I),
    .ce(CE),
    .out(value__CE_out),
    .clk(CLK)
);
assign O = value__CE_out;
endmodule

module RMUX_T4_WEST_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[19];
endmodule

module RMUX_T4_WEST_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[19];
endmodule

module RMUX_T4_SOUTH_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[18];
endmodule

module RMUX_T4_SOUTH_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[18];
endmodule

module RMUX_T4_NORTH_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[17];
endmodule

module RMUX_T4_NORTH_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[17];
endmodule

module RMUX_T4_EAST_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[16];
endmodule

module RMUX_T4_EAST_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[16];
endmodule

module RMUX_T3_WEST_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[15];
endmodule

module RMUX_T3_WEST_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[15];
endmodule

module RMUX_T3_SOUTH_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[14];
endmodule

module RMUX_T3_SOUTH_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[14];
endmodule

module RMUX_T3_NORTH_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[13];
endmodule

module RMUX_T3_NORTH_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[13];
endmodule

module RMUX_T3_EAST_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[12];
endmodule

module RMUX_T3_EAST_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[12];
endmodule

module RMUX_T2_WEST_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[11];
endmodule

module RMUX_T2_WEST_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[11];
endmodule

module RMUX_T2_SOUTH_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[10];
endmodule

module RMUX_T2_SOUTH_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[10];
endmodule

module RMUX_T2_NORTH_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[9];
endmodule

module RMUX_T2_NORTH_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[9];
endmodule

module RMUX_T2_EAST_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[8];
endmodule

module RMUX_T2_EAST_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[8];
endmodule

module RMUX_T1_WEST_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[7];
endmodule

module RMUX_T1_WEST_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[7];
endmodule

module RMUX_T1_SOUTH_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[6];
endmodule

module RMUX_T1_SOUTH_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[6];
endmodule

module RMUX_T1_NORTH_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[5];
endmodule

module RMUX_T1_NORTH_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[5];
endmodule

module RMUX_T1_EAST_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[4];
endmodule

module RMUX_T1_EAST_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[4];
endmodule

module RMUX_T0_WEST_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[3];
endmodule

module RMUX_T0_WEST_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[3];
endmodule

module RMUX_T0_SOUTH_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[2];
endmodule

module RMUX_T0_SOUTH_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[2];
endmodule

module RMUX_T0_NORTH_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[1];
endmodule

module RMUX_T0_NORTH_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[1];
endmodule

module RMUX_T0_EAST_B1_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[0];
endmodule

module RMUX_T0_EAST_B16_sel (
    input [31:0] I,
    output [0:0] O
);
assign O = I[0];
endmodule

module Or3x8 (
    input [7:0] I0,
    input [7:0] I1,
    input [7:0] I2,
    output [7:0] O
);
wire orr_inst0_out;
wire orr_inst1_out;
wire orr_inst2_out;
wire orr_inst3_out;
wire orr_inst4_out;
wire orr_inst5_out;
wire orr_inst6_out;
wire orr_inst7_out;
wire [2:0] orr_inst0_in;
assign orr_inst0_in = {I2[0],I1[0],I0[0]};
coreir_orr #(
    .width(3)
) orr_inst0 (
    .in(orr_inst0_in),
    .out(orr_inst0_out)
);
wire [2:0] orr_inst1_in;
assign orr_inst1_in = {I2[1],I1[1],I0[1]};
coreir_orr #(
    .width(3)
) orr_inst1 (
    .in(orr_inst1_in),
    .out(orr_inst1_out)
);
wire [2:0] orr_inst2_in;
assign orr_inst2_in = {I2[2],I1[2],I0[2]};
coreir_orr #(
    .width(3)
) orr_inst2 (
    .in(orr_inst2_in),
    .out(orr_inst2_out)
);
wire [2:0] orr_inst3_in;
assign orr_inst3_in = {I2[3],I1[3],I0[3]};
coreir_orr #(
    .width(3)
) orr_inst3 (
    .in(orr_inst3_in),
    .out(orr_inst3_out)
);
wire [2:0] orr_inst4_in;
assign orr_inst4_in = {I2[4],I1[4],I0[4]};
coreir_orr #(
    .width(3)
) orr_inst4 (
    .in(orr_inst4_in),
    .out(orr_inst4_out)
);
wire [2:0] orr_inst5_in;
assign orr_inst5_in = {I2[5],I1[5],I0[5]};
coreir_orr #(
    .width(3)
) orr_inst5 (
    .in(orr_inst5_in),
    .out(orr_inst5_out)
);
wire [2:0] orr_inst6_in;
assign orr_inst6_in = {I2[6],I1[6],I0[6]};
coreir_orr #(
    .width(3)
) orr_inst6 (
    .in(orr_inst6_in),
    .out(orr_inst6_out)
);
wire [2:0] orr_inst7_in;
assign orr_inst7_in = {I2[7],I1[7],I0[7]};
coreir_orr #(
    .width(3)
) orr_inst7 (
    .in(orr_inst7_in),
    .out(orr_inst7_out)
);
assign O = {orr_inst7_out,orr_inst6_out,orr_inst5_out,orr_inst4_out,orr_inst3_out,orr_inst2_out,orr_inst1_out,orr_inst0_out};
endmodule

module Or3x32 (
    input [31:0] I0,
    input [31:0] I1,
    input [31:0] I2,
    output [31:0] O
);
wire orr_inst0_out;
wire orr_inst1_out;
wire orr_inst10_out;
wire orr_inst11_out;
wire orr_inst12_out;
wire orr_inst13_out;
wire orr_inst14_out;
wire orr_inst15_out;
wire orr_inst16_out;
wire orr_inst17_out;
wire orr_inst18_out;
wire orr_inst19_out;
wire orr_inst2_out;
wire orr_inst20_out;
wire orr_inst21_out;
wire orr_inst22_out;
wire orr_inst23_out;
wire orr_inst24_out;
wire orr_inst25_out;
wire orr_inst26_out;
wire orr_inst27_out;
wire orr_inst28_out;
wire orr_inst29_out;
wire orr_inst3_out;
wire orr_inst30_out;
wire orr_inst31_out;
wire orr_inst4_out;
wire orr_inst5_out;
wire orr_inst6_out;
wire orr_inst7_out;
wire orr_inst8_out;
wire orr_inst9_out;
wire [2:0] orr_inst0_in;
assign orr_inst0_in = {I2[0],I1[0],I0[0]};
coreir_orr #(
    .width(3)
) orr_inst0 (
    .in(orr_inst0_in),
    .out(orr_inst0_out)
);
wire [2:0] orr_inst1_in;
assign orr_inst1_in = {I2[1],I1[1],I0[1]};
coreir_orr #(
    .width(3)
) orr_inst1 (
    .in(orr_inst1_in),
    .out(orr_inst1_out)
);
wire [2:0] orr_inst10_in;
assign orr_inst10_in = {I2[10],I1[10],I0[10]};
coreir_orr #(
    .width(3)
) orr_inst10 (
    .in(orr_inst10_in),
    .out(orr_inst10_out)
);
wire [2:0] orr_inst11_in;
assign orr_inst11_in = {I2[11],I1[11],I0[11]};
coreir_orr #(
    .width(3)
) orr_inst11 (
    .in(orr_inst11_in),
    .out(orr_inst11_out)
);
wire [2:0] orr_inst12_in;
assign orr_inst12_in = {I2[12],I1[12],I0[12]};
coreir_orr #(
    .width(3)
) orr_inst12 (
    .in(orr_inst12_in),
    .out(orr_inst12_out)
);
wire [2:0] orr_inst13_in;
assign orr_inst13_in = {I2[13],I1[13],I0[13]};
coreir_orr #(
    .width(3)
) orr_inst13 (
    .in(orr_inst13_in),
    .out(orr_inst13_out)
);
wire [2:0] orr_inst14_in;
assign orr_inst14_in = {I2[14],I1[14],I0[14]};
coreir_orr #(
    .width(3)
) orr_inst14 (
    .in(orr_inst14_in),
    .out(orr_inst14_out)
);
wire [2:0] orr_inst15_in;
assign orr_inst15_in = {I2[15],I1[15],I0[15]};
coreir_orr #(
    .width(3)
) orr_inst15 (
    .in(orr_inst15_in),
    .out(orr_inst15_out)
);
wire [2:0] orr_inst16_in;
assign orr_inst16_in = {I2[16],I1[16],I0[16]};
coreir_orr #(
    .width(3)
) orr_inst16 (
    .in(orr_inst16_in),
    .out(orr_inst16_out)
);
wire [2:0] orr_inst17_in;
assign orr_inst17_in = {I2[17],I1[17],I0[17]};
coreir_orr #(
    .width(3)
) orr_inst17 (
    .in(orr_inst17_in),
    .out(orr_inst17_out)
);
wire [2:0] orr_inst18_in;
assign orr_inst18_in = {I2[18],I1[18],I0[18]};
coreir_orr #(
    .width(3)
) orr_inst18 (
    .in(orr_inst18_in),
    .out(orr_inst18_out)
);
wire [2:0] orr_inst19_in;
assign orr_inst19_in = {I2[19],I1[19],I0[19]};
coreir_orr #(
    .width(3)
) orr_inst19 (
    .in(orr_inst19_in),
    .out(orr_inst19_out)
);
wire [2:0] orr_inst2_in;
assign orr_inst2_in = {I2[2],I1[2],I0[2]};
coreir_orr #(
    .width(3)
) orr_inst2 (
    .in(orr_inst2_in),
    .out(orr_inst2_out)
);
wire [2:0] orr_inst20_in;
assign orr_inst20_in = {I2[20],I1[20],I0[20]};
coreir_orr #(
    .width(3)
) orr_inst20 (
    .in(orr_inst20_in),
    .out(orr_inst20_out)
);
wire [2:0] orr_inst21_in;
assign orr_inst21_in = {I2[21],I1[21],I0[21]};
coreir_orr #(
    .width(3)
) orr_inst21 (
    .in(orr_inst21_in),
    .out(orr_inst21_out)
);
wire [2:0] orr_inst22_in;
assign orr_inst22_in = {I2[22],I1[22],I0[22]};
coreir_orr #(
    .width(3)
) orr_inst22 (
    .in(orr_inst22_in),
    .out(orr_inst22_out)
);
wire [2:0] orr_inst23_in;
assign orr_inst23_in = {I2[23],I1[23],I0[23]};
coreir_orr #(
    .width(3)
) orr_inst23 (
    .in(orr_inst23_in),
    .out(orr_inst23_out)
);
wire [2:0] orr_inst24_in;
assign orr_inst24_in = {I2[24],I1[24],I0[24]};
coreir_orr #(
    .width(3)
) orr_inst24 (
    .in(orr_inst24_in),
    .out(orr_inst24_out)
);
wire [2:0] orr_inst25_in;
assign orr_inst25_in = {I2[25],I1[25],I0[25]};
coreir_orr #(
    .width(3)
) orr_inst25 (
    .in(orr_inst25_in),
    .out(orr_inst25_out)
);
wire [2:0] orr_inst26_in;
assign orr_inst26_in = {I2[26],I1[26],I0[26]};
coreir_orr #(
    .width(3)
) orr_inst26 (
    .in(orr_inst26_in),
    .out(orr_inst26_out)
);
wire [2:0] orr_inst27_in;
assign orr_inst27_in = {I2[27],I1[27],I0[27]};
coreir_orr #(
    .width(3)
) orr_inst27 (
    .in(orr_inst27_in),
    .out(orr_inst27_out)
);
wire [2:0] orr_inst28_in;
assign orr_inst28_in = {I2[28],I1[28],I0[28]};
coreir_orr #(
    .width(3)
) orr_inst28 (
    .in(orr_inst28_in),
    .out(orr_inst28_out)
);
wire [2:0] orr_inst29_in;
assign orr_inst29_in = {I2[29],I1[29],I0[29]};
coreir_orr #(
    .width(3)
) orr_inst29 (
    .in(orr_inst29_in),
    .out(orr_inst29_out)
);
wire [2:0] orr_inst3_in;
assign orr_inst3_in = {I2[3],I1[3],I0[3]};
coreir_orr #(
    .width(3)
) orr_inst3 (
    .in(orr_inst3_in),
    .out(orr_inst3_out)
);
wire [2:0] orr_inst30_in;
assign orr_inst30_in = {I2[30],I1[30],I0[30]};
coreir_orr #(
    .width(3)
) orr_inst30 (
    .in(orr_inst30_in),
    .out(orr_inst30_out)
);
wire [2:0] orr_inst31_in;
assign orr_inst31_in = {I2[31],I1[31],I0[31]};
coreir_orr #(
    .width(3)
) orr_inst31 (
    .in(orr_inst31_in),
    .out(orr_inst31_out)
);
wire [2:0] orr_inst4_in;
assign orr_inst4_in = {I2[4],I1[4],I0[4]};
coreir_orr #(
    .width(3)
) orr_inst4 (
    .in(orr_inst4_in),
    .out(orr_inst4_out)
);
wire [2:0] orr_inst5_in;
assign orr_inst5_in = {I2[5],I1[5],I0[5]};
coreir_orr #(
    .width(3)
) orr_inst5 (
    .in(orr_inst5_in),
    .out(orr_inst5_out)
);
wire [2:0] orr_inst6_in;
assign orr_inst6_in = {I2[6],I1[6],I0[6]};
coreir_orr #(
    .width(3)
) orr_inst6 (
    .in(orr_inst6_in),
    .out(orr_inst6_out)
);
wire [2:0] orr_inst7_in;
assign orr_inst7_in = {I2[7],I1[7],I0[7]};
coreir_orr #(
    .width(3)
) orr_inst7 (
    .in(orr_inst7_in),
    .out(orr_inst7_out)
);
wire [2:0] orr_inst8_in;
assign orr_inst8_in = {I2[8],I1[8],I0[8]};
coreir_orr #(
    .width(3)
) orr_inst8 (
    .in(orr_inst8_in),
    .out(orr_inst8_out)
);
wire [2:0] orr_inst9_in;
assign orr_inst9_in = {I2[9],I1[9],I0[9]};
coreir_orr #(
    .width(3)
) orr_inst9 (
    .in(orr_inst9_in),
    .out(orr_inst9_out)
);
assign O = {orr_inst31_out,orr_inst30_out,orr_inst29_out,orr_inst28_out,orr_inst27_out,orr_inst26_out,orr_inst25_out,orr_inst24_out,orr_inst23_out,orr_inst22_out,orr_inst21_out,orr_inst20_out,orr_inst19_out,orr_inst18_out,orr_inst17_out,orr_inst16_out,orr_inst15_out,orr_inst14_out,orr_inst13_out,orr_inst12_out,orr_inst11_out,orr_inst10_out,orr_inst9_out,orr_inst8_out,orr_inst7_out,orr_inst6_out,orr_inst5_out,orr_inst4_out,orr_inst3_out,orr_inst2_out,orr_inst1_out,orr_inst0_out};
endmodule

module Or16x32 (
    input [31:0] I0,
    input [31:0] I1,
    input [31:0] I2,
    input [31:0] I3,
    input [31:0] I4,
    input [31:0] I5,
    input [31:0] I6,
    input [31:0] I7,
    input [31:0] I8,
    input [31:0] I9,
    input [31:0] I10,
    input [31:0] I11,
    input [31:0] I12,
    input [31:0] I13,
    input [31:0] I14,
    input [31:0] I15,
    output [31:0] O
);
wire orr_inst0_out;
wire orr_inst1_out;
wire orr_inst10_out;
wire orr_inst11_out;
wire orr_inst12_out;
wire orr_inst13_out;
wire orr_inst14_out;
wire orr_inst15_out;
wire orr_inst16_out;
wire orr_inst17_out;
wire orr_inst18_out;
wire orr_inst19_out;
wire orr_inst2_out;
wire orr_inst20_out;
wire orr_inst21_out;
wire orr_inst22_out;
wire orr_inst23_out;
wire orr_inst24_out;
wire orr_inst25_out;
wire orr_inst26_out;
wire orr_inst27_out;
wire orr_inst28_out;
wire orr_inst29_out;
wire orr_inst3_out;
wire orr_inst30_out;
wire orr_inst31_out;
wire orr_inst4_out;
wire orr_inst5_out;
wire orr_inst6_out;
wire orr_inst7_out;
wire orr_inst8_out;
wire orr_inst9_out;
wire [15:0] orr_inst0_in;
assign orr_inst0_in = {I15[0],I14[0],I13[0],I12[0],I11[0],I10[0],I9[0],I8[0],I7[0],I6[0],I5[0],I4[0],I3[0],I2[0],I1[0],I0[0]};
coreir_orr #(
    .width(16)
) orr_inst0 (
    .in(orr_inst0_in),
    .out(orr_inst0_out)
);
wire [15:0] orr_inst1_in;
assign orr_inst1_in = {I15[1],I14[1],I13[1],I12[1],I11[1],I10[1],I9[1],I8[1],I7[1],I6[1],I5[1],I4[1],I3[1],I2[1],I1[1],I0[1]};
coreir_orr #(
    .width(16)
) orr_inst1 (
    .in(orr_inst1_in),
    .out(orr_inst1_out)
);
wire [15:0] orr_inst10_in;
assign orr_inst10_in = {I15[10],I14[10],I13[10],I12[10],I11[10],I10[10],I9[10],I8[10],I7[10],I6[10],I5[10],I4[10],I3[10],I2[10],I1[10],I0[10]};
coreir_orr #(
    .width(16)
) orr_inst10 (
    .in(orr_inst10_in),
    .out(orr_inst10_out)
);
wire [15:0] orr_inst11_in;
assign orr_inst11_in = {I15[11],I14[11],I13[11],I12[11],I11[11],I10[11],I9[11],I8[11],I7[11],I6[11],I5[11],I4[11],I3[11],I2[11],I1[11],I0[11]};
coreir_orr #(
    .width(16)
) orr_inst11 (
    .in(orr_inst11_in),
    .out(orr_inst11_out)
);
wire [15:0] orr_inst12_in;
assign orr_inst12_in = {I15[12],I14[12],I13[12],I12[12],I11[12],I10[12],I9[12],I8[12],I7[12],I6[12],I5[12],I4[12],I3[12],I2[12],I1[12],I0[12]};
coreir_orr #(
    .width(16)
) orr_inst12 (
    .in(orr_inst12_in),
    .out(orr_inst12_out)
);
wire [15:0] orr_inst13_in;
assign orr_inst13_in = {I15[13],I14[13],I13[13],I12[13],I11[13],I10[13],I9[13],I8[13],I7[13],I6[13],I5[13],I4[13],I3[13],I2[13],I1[13],I0[13]};
coreir_orr #(
    .width(16)
) orr_inst13 (
    .in(orr_inst13_in),
    .out(orr_inst13_out)
);
wire [15:0] orr_inst14_in;
assign orr_inst14_in = {I15[14],I14[14],I13[14],I12[14],I11[14],I10[14],I9[14],I8[14],I7[14],I6[14],I5[14],I4[14],I3[14],I2[14],I1[14],I0[14]};
coreir_orr #(
    .width(16)
) orr_inst14 (
    .in(orr_inst14_in),
    .out(orr_inst14_out)
);
wire [15:0] orr_inst15_in;
assign orr_inst15_in = {I15[15],I14[15],I13[15],I12[15],I11[15],I10[15],I9[15],I8[15],I7[15],I6[15],I5[15],I4[15],I3[15],I2[15],I1[15],I0[15]};
coreir_orr #(
    .width(16)
) orr_inst15 (
    .in(orr_inst15_in),
    .out(orr_inst15_out)
);
wire [15:0] orr_inst16_in;
assign orr_inst16_in = {I15[16],I14[16],I13[16],I12[16],I11[16],I10[16],I9[16],I8[16],I7[16],I6[16],I5[16],I4[16],I3[16],I2[16],I1[16],I0[16]};
coreir_orr #(
    .width(16)
) orr_inst16 (
    .in(orr_inst16_in),
    .out(orr_inst16_out)
);
wire [15:0] orr_inst17_in;
assign orr_inst17_in = {I15[17],I14[17],I13[17],I12[17],I11[17],I10[17],I9[17],I8[17],I7[17],I6[17],I5[17],I4[17],I3[17],I2[17],I1[17],I0[17]};
coreir_orr #(
    .width(16)
) orr_inst17 (
    .in(orr_inst17_in),
    .out(orr_inst17_out)
);
wire [15:0] orr_inst18_in;
assign orr_inst18_in = {I15[18],I14[18],I13[18],I12[18],I11[18],I10[18],I9[18],I8[18],I7[18],I6[18],I5[18],I4[18],I3[18],I2[18],I1[18],I0[18]};
coreir_orr #(
    .width(16)
) orr_inst18 (
    .in(orr_inst18_in),
    .out(orr_inst18_out)
);
wire [15:0] orr_inst19_in;
assign orr_inst19_in = {I15[19],I14[19],I13[19],I12[19],I11[19],I10[19],I9[19],I8[19],I7[19],I6[19],I5[19],I4[19],I3[19],I2[19],I1[19],I0[19]};
coreir_orr #(
    .width(16)
) orr_inst19 (
    .in(orr_inst19_in),
    .out(orr_inst19_out)
);
wire [15:0] orr_inst2_in;
assign orr_inst2_in = {I15[2],I14[2],I13[2],I12[2],I11[2],I10[2],I9[2],I8[2],I7[2],I6[2],I5[2],I4[2],I3[2],I2[2],I1[2],I0[2]};
coreir_orr #(
    .width(16)
) orr_inst2 (
    .in(orr_inst2_in),
    .out(orr_inst2_out)
);
wire [15:0] orr_inst20_in;
assign orr_inst20_in = {I15[20],I14[20],I13[20],I12[20],I11[20],I10[20],I9[20],I8[20],I7[20],I6[20],I5[20],I4[20],I3[20],I2[20],I1[20],I0[20]};
coreir_orr #(
    .width(16)
) orr_inst20 (
    .in(orr_inst20_in),
    .out(orr_inst20_out)
);
wire [15:0] orr_inst21_in;
assign orr_inst21_in = {I15[21],I14[21],I13[21],I12[21],I11[21],I10[21],I9[21],I8[21],I7[21],I6[21],I5[21],I4[21],I3[21],I2[21],I1[21],I0[21]};
coreir_orr #(
    .width(16)
) orr_inst21 (
    .in(orr_inst21_in),
    .out(orr_inst21_out)
);
wire [15:0] orr_inst22_in;
assign orr_inst22_in = {I15[22],I14[22],I13[22],I12[22],I11[22],I10[22],I9[22],I8[22],I7[22],I6[22],I5[22],I4[22],I3[22],I2[22],I1[22],I0[22]};
coreir_orr #(
    .width(16)
) orr_inst22 (
    .in(orr_inst22_in),
    .out(orr_inst22_out)
);
wire [15:0] orr_inst23_in;
assign orr_inst23_in = {I15[23],I14[23],I13[23],I12[23],I11[23],I10[23],I9[23],I8[23],I7[23],I6[23],I5[23],I4[23],I3[23],I2[23],I1[23],I0[23]};
coreir_orr #(
    .width(16)
) orr_inst23 (
    .in(orr_inst23_in),
    .out(orr_inst23_out)
);
wire [15:0] orr_inst24_in;
assign orr_inst24_in = {I15[24],I14[24],I13[24],I12[24],I11[24],I10[24],I9[24],I8[24],I7[24],I6[24],I5[24],I4[24],I3[24],I2[24],I1[24],I0[24]};
coreir_orr #(
    .width(16)
) orr_inst24 (
    .in(orr_inst24_in),
    .out(orr_inst24_out)
);
wire [15:0] orr_inst25_in;
assign orr_inst25_in = {I15[25],I14[25],I13[25],I12[25],I11[25],I10[25],I9[25],I8[25],I7[25],I6[25],I5[25],I4[25],I3[25],I2[25],I1[25],I0[25]};
coreir_orr #(
    .width(16)
) orr_inst25 (
    .in(orr_inst25_in),
    .out(orr_inst25_out)
);
wire [15:0] orr_inst26_in;
assign orr_inst26_in = {I15[26],I14[26],I13[26],I12[26],I11[26],I10[26],I9[26],I8[26],I7[26],I6[26],I5[26],I4[26],I3[26],I2[26],I1[26],I0[26]};
coreir_orr #(
    .width(16)
) orr_inst26 (
    .in(orr_inst26_in),
    .out(orr_inst26_out)
);
wire [15:0] orr_inst27_in;
assign orr_inst27_in = {I15[27],I14[27],I13[27],I12[27],I11[27],I10[27],I9[27],I8[27],I7[27],I6[27],I5[27],I4[27],I3[27],I2[27],I1[27],I0[27]};
coreir_orr #(
    .width(16)
) orr_inst27 (
    .in(orr_inst27_in),
    .out(orr_inst27_out)
);
wire [15:0] orr_inst28_in;
assign orr_inst28_in = {I15[28],I14[28],I13[28],I12[28],I11[28],I10[28],I9[28],I8[28],I7[28],I6[28],I5[28],I4[28],I3[28],I2[28],I1[28],I0[28]};
coreir_orr #(
    .width(16)
) orr_inst28 (
    .in(orr_inst28_in),
    .out(orr_inst28_out)
);
wire [15:0] orr_inst29_in;
assign orr_inst29_in = {I15[29],I14[29],I13[29],I12[29],I11[29],I10[29],I9[29],I8[29],I7[29],I6[29],I5[29],I4[29],I3[29],I2[29],I1[29],I0[29]};
coreir_orr #(
    .width(16)
) orr_inst29 (
    .in(orr_inst29_in),
    .out(orr_inst29_out)
);
wire [15:0] orr_inst3_in;
assign orr_inst3_in = {I15[3],I14[3],I13[3],I12[3],I11[3],I10[3],I9[3],I8[3],I7[3],I6[3],I5[3],I4[3],I3[3],I2[3],I1[3],I0[3]};
coreir_orr #(
    .width(16)
) orr_inst3 (
    .in(orr_inst3_in),
    .out(orr_inst3_out)
);
wire [15:0] orr_inst30_in;
assign orr_inst30_in = {I15[30],I14[30],I13[30],I12[30],I11[30],I10[30],I9[30],I8[30],I7[30],I6[30],I5[30],I4[30],I3[30],I2[30],I1[30],I0[30]};
coreir_orr #(
    .width(16)
) orr_inst30 (
    .in(orr_inst30_in),
    .out(orr_inst30_out)
);
wire [15:0] orr_inst31_in;
assign orr_inst31_in = {I15[31],I14[31],I13[31],I12[31],I11[31],I10[31],I9[31],I8[31],I7[31],I6[31],I5[31],I4[31],I3[31],I2[31],I1[31],I0[31]};
coreir_orr #(
    .width(16)
) orr_inst31 (
    .in(orr_inst31_in),
    .out(orr_inst31_out)
);
wire [15:0] orr_inst4_in;
assign orr_inst4_in = {I15[4],I14[4],I13[4],I12[4],I11[4],I10[4],I9[4],I8[4],I7[4],I6[4],I5[4],I4[4],I3[4],I2[4],I1[4],I0[4]};
coreir_orr #(
    .width(16)
) orr_inst4 (
    .in(orr_inst4_in),
    .out(orr_inst4_out)
);
wire [15:0] orr_inst5_in;
assign orr_inst5_in = {I15[5],I14[5],I13[5],I12[5],I11[5],I10[5],I9[5],I8[5],I7[5],I6[5],I5[5],I4[5],I3[5],I2[5],I1[5],I0[5]};
coreir_orr #(
    .width(16)
) orr_inst5 (
    .in(orr_inst5_in),
    .out(orr_inst5_out)
);
wire [15:0] orr_inst6_in;
assign orr_inst6_in = {I15[6],I14[6],I13[6],I12[6],I11[6],I10[6],I9[6],I8[6],I7[6],I6[6],I5[6],I4[6],I3[6],I2[6],I1[6],I0[6]};
coreir_orr #(
    .width(16)
) orr_inst6 (
    .in(orr_inst6_in),
    .out(orr_inst6_out)
);
wire [15:0] orr_inst7_in;
assign orr_inst7_in = {I15[7],I14[7],I13[7],I12[7],I11[7],I10[7],I9[7],I8[7],I7[7],I6[7],I5[7],I4[7],I3[7],I2[7],I1[7],I0[7]};
coreir_orr #(
    .width(16)
) orr_inst7 (
    .in(orr_inst7_in),
    .out(orr_inst7_out)
);
wire [15:0] orr_inst8_in;
assign orr_inst8_in = {I15[8],I14[8],I13[8],I12[8],I11[8],I10[8],I9[8],I8[8],I7[8],I6[8],I5[8],I4[8],I3[8],I2[8],I1[8],I0[8]};
coreir_orr #(
    .width(16)
) orr_inst8 (
    .in(orr_inst8_in),
    .out(orr_inst8_out)
);
wire [15:0] orr_inst9_in;
assign orr_inst9_in = {I15[9],I14[9],I13[9],I12[9],I11[9],I10[9],I9[9],I8[9],I7[9],I6[9],I5[9],I4[9],I3[9],I2[9],I1[9],I0[9]};
coreir_orr #(
    .width(16)
) orr_inst9 (
    .in(orr_inst9_in),
    .out(orr_inst9_out)
);
assign O = {orr_inst31_out,orr_inst30_out,orr_inst29_out,orr_inst28_out,orr_inst27_out,orr_inst26_out,orr_inst25_out,orr_inst24_out,orr_inst23_out,orr_inst22_out,orr_inst21_out,orr_inst20_out,orr_inst19_out,orr_inst18_out,orr_inst17_out,orr_inst16_out,orr_inst15_out,orr_inst14_out,orr_inst13_out,orr_inst12_out,orr_inst11_out,orr_inst10_out,orr_inst9_out,orr_inst8_out,orr_inst7_out,orr_inst6_out,orr_inst5_out,orr_inst4_out,orr_inst3_out,orr_inst2_out,orr_inst1_out,orr_inst0_out};
endmodule

module MuxWrapper_1_16 (
    input [15:0] I,
    output [15:0] O
);
assign O = I;
endmodule

module MuxWrapper_1_1 (
    input [0:0] I,
    output [0:0] O
);
assign O = I;
endmodule

module Tile_io_core (
    input [15:0] tile_id,
    input [0:0] glb2io_1,
    input [0:0] f2io_1,
    output [0:0] io2glb_1,
    output [0:0] io2f_1,
    input [15:0] glb2io_16,
    input [15:0] f2io_16,
    output [15:0] io2glb_16,
    output [15:0] io2f_16,
    output [8:0] hi,
    output [7:0] lo
);
wire [0:0] CB_f2io_1$WIRE_CB_f2io_1_O;
wire [15:0] CB_f2io_16$WIRE_CB_f2io_16_O;
wire [7:0] const_0_8_out;
wire [8:0] const_511_9_out;
wire [15:0] io_core_inst0_io2glb_16;
wire [0:0] io_core_inst0_io2glb_1;
wire [15:0] io_core_inst0_io2f_16;
wire [0:0] io_core_inst0_io2f_1;
MuxWrapper_1_1 CB_f2io_1$WIRE_CB_f2io_1 (
    .I(f2io_1),
    .O(CB_f2io_1$WIRE_CB_f2io_1_O)
);
MuxWrapper_1_16 CB_f2io_16$WIRE_CB_f2io_16 (
    .I(f2io_16),
    .O(CB_f2io_16$WIRE_CB_f2io_16_O)
);
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
coreir_const #(
    .value(9'h1ff),
    .width(9)
) const_511_9 (
    .out(const_511_9_out)
);
io_core io_core_inst0 (
    .glb2io_16(glb2io_16),
    .glb2io_1(glb2io_1),
    .io2glb_16(io_core_inst0_io2glb_16),
    .io2glb_1(io_core_inst0_io2glb_1),
    .f2io_16(CB_f2io_16$WIRE_CB_f2io_16_O),
    .f2io_1(CB_f2io_1$WIRE_CB_f2io_1_O),
    .io2f_16(io_core_inst0_io2f_16),
    .io2f_1(io_core_inst0_io2f_1)
);
assign io2glb_1 = io_core_inst0_io2glb_1;
assign io2f_1 = io_core_inst0_io2f_1;
assign io2glb_16 = io_core_inst0_io2glb_16;
assign io2f_16 = io_core_inst0_io2f_16;
assign hi = const_511_9_out;
assign lo = const_0_8_out;
endmodule

module MuxWithDefaultWrapper_9_32_8_0 (
    input [0:0] EN,
    input [31:0] I_0,
    input [31:0] I_1,
    input [31:0] I_2,
    input [31:0] I_3,
    input [31:0] I_4,
    input [31:0] I_5,
    input [31:0] I_6,
    input [31:0] I_7,
    input [31:0] I_8,
    output [31:0] O,
    input [7:0] S
);
wire [31:0] MuxWrapper_2_32_inst0$Mux2x32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
wire [31:0] MuxWrapper_9_32_inst0$Mux9x32_inst0$coreir_commonlib_mux9x32_inst0_out;
wire [3:0] MuxWrapper_9_32_inst0_S_in;
wire and_inst0_out;
wire [31:0] const_0_32_out;
wire [7:0] const_9_8_out;
wire coreir_ult8_inst0_out;
wire [7:0] self_S_out;
coreir_mux #(
    .width(32)
) MuxWrapper_2_32_inst0$Mux2x32_inst0$coreir_commonlib_mux2x32_inst0$_join (
    .in0(const_0_32_out),
    .in1(MuxWrapper_9_32_inst0$Mux9x32_inst0$coreir_commonlib_mux9x32_inst0_out),
    .sel(and_inst0_out),
    .out(MuxWrapper_2_32_inst0$Mux2x32_inst0$coreir_commonlib_mux2x32_inst0$_join_out)
);
commonlib_muxn__N9__width32 MuxWrapper_9_32_inst0$Mux9x32_inst0$coreir_commonlib_mux9x32_inst0 (
    .in_data_0(I_0),
    .in_data_1(I_1),
    .in_data_2(I_2),
    .in_data_3(I_3),
    .in_data_4(I_4),
    .in_data_5(I_5),
    .in_data_6(I_6),
    .in_data_7(I_7),
    .in_data_8(I_8),
    .in_sel(MuxWrapper_9_32_inst0_S_in),
    .out(MuxWrapper_9_32_inst0$Mux9x32_inst0$coreir_commonlib_mux9x32_inst0_out)
);
mantle_wire__typeBitIn4 MuxWrapper_9_32_inst0_S (
    .in(MuxWrapper_9_32_inst0_S_in),
    .out(self_S_out[3:0])
);
corebit_and and_inst0 (
    .in0(coreir_ult8_inst0_out),
    .in1(EN[0]),
    .out(and_inst0_out)
);
coreir_const #(
    .value(32'h00000000),
    .width(32)
) const_0_32 (
    .out(const_0_32_out)
);
coreir_const #(
    .value(8'h09),
    .width(8)
) const_9_8 (
    .out(const_9_8_out)
);
coreir_ult #(
    .width(8)
) coreir_ult8_inst0 (
    .in0(S),
    .in1(const_9_8_out),
    .out(coreir_ult8_inst0_out)
);
mantle_wire__typeBit8 self_S (
    .in(S),
    .out(self_S_out)
);
assign O = MuxWrapper_2_32_inst0$Mux2x32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
endmodule

module MuxWithDefaultWrapper_16_32_8_0 (
    input [0:0] EN,
    input [31:0] I_0,
    input [31:0] I_1,
    input [31:0] I_10,
    input [31:0] I_11,
    input [31:0] I_12,
    input [31:0] I_13,
    input [31:0] I_14,
    input [31:0] I_15,
    input [31:0] I_2,
    input [31:0] I_3,
    input [31:0] I_4,
    input [31:0] I_5,
    input [31:0] I_6,
    input [31:0] I_7,
    input [31:0] I_8,
    input [31:0] I_9,
    output [31:0] O,
    input [7:0] S
);
wire [31:0] MuxWrapper_16_32_inst0$Mux16x32_inst0$coreir_commonlib_mux16x32_inst0_out;
wire [3:0] MuxWrapper_16_32_inst0_S_in;
wire [31:0] MuxWrapper_2_32_inst0$Mux2x32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
wire and_inst0_out;
wire [31:0] const_0_32_out;
wire [7:0] const_16_8_out;
wire coreir_ult8_inst0_out;
wire [7:0] self_S_out;
commonlib_muxn__N16__width32 MuxWrapper_16_32_inst0$Mux16x32_inst0$coreir_commonlib_mux16x32_inst0 (
    .in_data_0(I_0),
    .in_data_1(I_1),
    .in_data_10(I_10),
    .in_data_11(I_11),
    .in_data_12(I_12),
    .in_data_13(I_13),
    .in_data_14(I_14),
    .in_data_15(I_15),
    .in_data_2(I_2),
    .in_data_3(I_3),
    .in_data_4(I_4),
    .in_data_5(I_5),
    .in_data_6(I_6),
    .in_data_7(I_7),
    .in_data_8(I_8),
    .in_data_9(I_9),
    .in_sel(MuxWrapper_16_32_inst0_S_in),
    .out(MuxWrapper_16_32_inst0$Mux16x32_inst0$coreir_commonlib_mux16x32_inst0_out)
);
mantle_wire__typeBitIn4 MuxWrapper_16_32_inst0_S (
    .in(MuxWrapper_16_32_inst0_S_in),
    .out(self_S_out[3:0])
);
coreir_mux #(
    .width(32)
) MuxWrapper_2_32_inst0$Mux2x32_inst0$coreir_commonlib_mux2x32_inst0$_join (
    .in0(const_0_32_out),
    .in1(MuxWrapper_16_32_inst0$Mux16x32_inst0$coreir_commonlib_mux16x32_inst0_out),
    .sel(and_inst0_out),
    .out(MuxWrapper_2_32_inst0$Mux2x32_inst0$coreir_commonlib_mux2x32_inst0$_join_out)
);
corebit_and and_inst0 (
    .in0(coreir_ult8_inst0_out),
    .in1(EN[0]),
    .out(and_inst0_out)
);
coreir_const #(
    .value(32'h00000000),
    .width(32)
) const_0_32 (
    .out(const_0_32_out)
);
coreir_const #(
    .value(8'h10),
    .width(8)
) const_16_8 (
    .out(const_16_8_out)
);
coreir_ult #(
    .width(8)
) coreir_ult8_inst0 (
    .in0(S),
    .in1(const_16_8_out),
    .out(coreir_ult8_inst0_out)
);
mantle_wire__typeBit8 self_S (
    .in(S),
    .out(self_S_out)
);
assign O = MuxWrapper_2_32_inst0$Mux2x32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
endmodule

module MUL (
    input [1:0] instr,
    input [0:0] signed_,
    input [15:0] a,
    input [15:0] b,
    output [15:0] O,
    input CLK,
    input ASYNCRESET
);
wire [15:0] Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst0_O_out;
wire [15:0] Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst1_O_out;
wire [15:0] Mux2xUInt16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xUInt16_inst0_I0_in;
wire [15:0] Mux2xUInt16_inst0_I1_in;
wire [31:0] Mux2xUInt32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
wire [31:0] Mux2xUInt32_inst0_I0_in;
wire [31:0] Mux2xUInt32_inst0_I1_in;
wire [31:0] Mux2xUInt32_inst1$coreir_commonlib_mux2x32_inst0$_join_out;
wire [31:0] Mux2xUInt32_inst1_I0_in;
wire [31:0] Mux2xUInt32_inst1_I1_in;
wire bit_const_0_None_out;
wire [15:0] const_0_16_out;
wire [1:0] const_0_2_out;
wire [0:0] const_1_1_out;
wire [1:0] const_2_2_out;
wire magma_Bits_1_eq_inst0_out;
wire magma_Bits_2_eq_inst0_out;
wire magma_Bits_2_eq_inst1_out;
wire [31:0] magma_Bits_32_and_inst0_out;
wire [31:0] magma_Bits_32_and_inst1_out;
wire [31:0] magma_Bits_32_mul_inst0_out;
coreir_mux #(
    .width(16)
) Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(a),
    .in1(const_0_16_out),
    .sel(magma_Bits_2_eq_inst0_out),
    .out(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
mantle_wire__typeBit16 Mux2xBits16_inst0_O (
    .in(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out),
    .out(Mux2xBits16_inst0_O_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join (
    .in0(b),
    .in1(const_0_16_out),
    .sel(magma_Bits_2_eq_inst0_out),
    .out(Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out)
);
mantle_wire__typeBit16 Mux2xBits16_inst1_O (
    .in(Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out),
    .out(Mux2xBits16_inst1_O_out)
);
coreir_mux #(
    .width(16)
) Mux2xUInt16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xUInt16_inst0_I0_in),
    .in1(Mux2xUInt16_inst0_I1_in),
    .sel(magma_Bits_2_eq_inst1_out),
    .out(Mux2xUInt16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
mantle_wire__typeBitIn16 Mux2xUInt16_inst0_I0 (
    .in(Mux2xUInt16_inst0_I0_in),
    .out(magma_Bits_32_mul_inst0_out[31:16])
);
mantle_wire__typeBitIn16 Mux2xUInt16_inst0_I1 (
    .in(Mux2xUInt16_inst0_I1_in),
    .out(magma_Bits_32_mul_inst0_out[15:0])
);
coreir_mux #(
    .width(32)
) Mux2xUInt32_inst0$coreir_commonlib_mux2x32_inst0$_join (
    .in0(Mux2xUInt32_inst0_I0_in),
    .in1(Mux2xUInt32_inst0_I1_in),
    .sel(magma_Bits_1_eq_inst0_out),
    .out(Mux2xUInt32_inst0$coreir_commonlib_mux2x32_inst0$_join_out)
);
wire [31:0] Mux2xUInt32_inst0_I0_out;
assign Mux2xUInt32_inst0_I0_out = {bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,Mux2xBits16_inst0_O_out[15:0]};
mantle_wire__typeBitIn32 Mux2xUInt32_inst0_I0 (
    .in(Mux2xUInt32_inst0_I0_in),
    .out(Mux2xUInt32_inst0_I0_out)
);
wire [31:0] Mux2xUInt32_inst0_I1_out;
assign Mux2xUInt32_inst0_I1_out = {Mux2xBits16_inst0_O_out[15],Mux2xBits16_inst0_O_out[15],Mux2xBits16_inst0_O_out[15],Mux2xBits16_inst0_O_out[15],Mux2xBits16_inst0_O_out[15],Mux2xBits16_inst0_O_out[15],Mux2xBits16_inst0_O_out[15],Mux2xBits16_inst0_O_out[15],Mux2xBits16_inst0_O_out[15],Mux2xBits16_inst0_O_out[15],Mux2xBits16_inst0_O_out[15],Mux2xBits16_inst0_O_out[15],Mux2xBits16_inst0_O_out[15],Mux2xBits16_inst0_O_out[15],Mux2xBits16_inst0_O_out[15],Mux2xBits16_inst0_O_out[15],Mux2xBits16_inst0_O_out[15:0]};
mantle_wire__typeBitIn32 Mux2xUInt32_inst0_I1 (
    .in(Mux2xUInt32_inst0_I1_in),
    .out(Mux2xUInt32_inst0_I1_out)
);
coreir_mux #(
    .width(32)
) Mux2xUInt32_inst1$coreir_commonlib_mux2x32_inst0$_join (
    .in0(Mux2xUInt32_inst1_I0_in),
    .in1(Mux2xUInt32_inst1_I1_in),
    .sel(magma_Bits_1_eq_inst0_out),
    .out(Mux2xUInt32_inst1$coreir_commonlib_mux2x32_inst0$_join_out)
);
wire [31:0] Mux2xUInt32_inst1_I0_out;
assign Mux2xUInt32_inst1_I0_out = {bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,Mux2xBits16_inst1_O_out[15:0]};
mantle_wire__typeBitIn32 Mux2xUInt32_inst1_I0 (
    .in(Mux2xUInt32_inst1_I0_in),
    .out(Mux2xUInt32_inst1_I0_out)
);
wire [31:0] Mux2xUInt32_inst1_I1_out;
assign Mux2xUInt32_inst1_I1_out = {Mux2xBits16_inst1_O_out[15],Mux2xBits16_inst1_O_out[15],Mux2xBits16_inst1_O_out[15],Mux2xBits16_inst1_O_out[15],Mux2xBits16_inst1_O_out[15],Mux2xBits16_inst1_O_out[15],Mux2xBits16_inst1_O_out[15],Mux2xBits16_inst1_O_out[15],Mux2xBits16_inst1_O_out[15],Mux2xBits16_inst1_O_out[15],Mux2xBits16_inst1_O_out[15],Mux2xBits16_inst1_O_out[15],Mux2xBits16_inst1_O_out[15],Mux2xBits16_inst1_O_out[15],Mux2xBits16_inst1_O_out[15],Mux2xBits16_inst1_O_out[15],Mux2xBits16_inst1_O_out[15:0]};
mantle_wire__typeBitIn32 Mux2xUInt32_inst1_I1 (
    .in(Mux2xUInt32_inst1_I1_in),
    .out(Mux2xUInt32_inst1_I1_out)
);
corebit_const #(
    .value(1'b0)
) bit_const_0_None (
    .out(bit_const_0_None_out)
);
coreir_const #(
    .value(16'h0000),
    .width(16)
) const_0_16 (
    .out(const_0_16_out)
);
coreir_const #(
    .value(2'h0),
    .width(2)
) const_0_2 (
    .out(const_0_2_out)
);
coreir_const #(
    .value(1'h1),
    .width(1)
) const_1_1 (
    .out(const_1_1_out)
);
coreir_const #(
    .value(2'h2),
    .width(2)
) const_2_2 (
    .out(const_2_2_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst0 (
    .in0(signed_),
    .in1(const_1_1_out),
    .out(magma_Bits_1_eq_inst0_out)
);
coreir_eq #(
    .width(2)
) magma_Bits_2_eq_inst0 (
    .in0(instr),
    .in1(const_2_2_out),
    .out(magma_Bits_2_eq_inst0_out)
);
coreir_eq #(
    .width(2)
) magma_Bits_2_eq_inst1 (
    .in0(instr),
    .in1(const_0_2_out),
    .out(magma_Bits_2_eq_inst1_out)
);
wire [31:0] magma_Bits_32_and_inst0_in1;
assign magma_Bits_32_and_inst0_in1 = {magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out};
coreir_and #(
    .width(32)
) magma_Bits_32_and_inst0 (
    .in0(Mux2xUInt32_inst0$coreir_commonlib_mux2x32_inst0$_join_out),
    .in1(magma_Bits_32_and_inst0_in1),
    .out(magma_Bits_32_and_inst0_out)
);
wire [31:0] magma_Bits_32_and_inst1_in1;
assign magma_Bits_32_and_inst1_in1 = {magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out,magma_Bits_2_eq_inst1_out};
coreir_and #(
    .width(32)
) magma_Bits_32_and_inst1 (
    .in0(Mux2xUInt32_inst1$coreir_commonlib_mux2x32_inst0$_join_out),
    .in1(magma_Bits_32_and_inst1_in1),
    .out(magma_Bits_32_and_inst1_out)
);
coreir_mul #(
    .width(32)
) magma_Bits_32_mul_inst0 (
    .in0(magma_Bits_32_and_inst0_out),
    .in1(magma_Bits_32_and_inst1_out),
    .out(magma_Bits_32_mul_inst0_out)
);
assign O = Mux2xUInt16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
endmodule

module Chain (
  input logic [1:0] accessor_output,
  input logic [1:0] [15:0] chain_data_in,
  input logic chain_en,
  input logic clk_en,
  input logic [1:0] [15:0] curr_tile_data_out,
  input logic flush,
  output logic [1:0] [15:0] data_out_tile
);

always_comb begin
  if (accessor_output[0]) begin
    data_out_tile[0] = curr_tile_data_out[0];
  end
  else if (chain_en) begin
    data_out_tile[0] = chain_data_in[0];
  end
  else data_out_tile[0] = 16'h0;
  if (accessor_output[1]) begin
    data_out_tile[1] = curr_tile_data_out[1];
  end
  else if (chain_en) begin
    data_out_tile[1] = chain_data_in[1];
  end
  else data_out_tile[1] = 16'h0;
end
endmodule   // Chain

module LakeTop (
  input logic [1:0] [15:0] addr_in,
  input logic chain_chain_en,
  input logic [1:0] [15:0] chain_data_in,
  input logic clk,
  input logic clk_en,
  input logic [7:0] config_addr_in,
  input logic [31:0] config_data_in,
  input logic [1:0] config_en,
  input logic config_read,
  input logic config_write,
  input logic [1:0] [15:0] data_in,
  input logic [15:0] fifo_ctrl_fifo_depth,
  input logic flush,
  input logic [3:0] loops_stencil_valid_dimensionality,
  input logic [5:0] [15:0] loops_stencil_valid_ranges,
  input logic [1:0] mode,
  input logic [1:0] ren_in,
  input logic rst_n,
  input logic stencil_valid_sched_gen_enable,
  input logic [15:0] stencil_valid_sched_gen_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] stencil_valid_sched_gen_sched_addr_gen_strides,
  input logic [3:0] strg_ub_agg_only_agg_read_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] strg_ub_agg_only_agg_read_addr_gen_0_strides,
  input logic [3:0] strg_ub_agg_only_agg_read_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] strg_ub_agg_only_agg_read_addr_gen_1_strides,
  input logic [3:0] strg_ub_agg_only_agg_write_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] strg_ub_agg_only_agg_write_addr_gen_0_strides,
  input logic [3:0] strg_ub_agg_only_agg_write_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] strg_ub_agg_only_agg_write_addr_gen_1_strides,
  input logic strg_ub_agg_only_agg_write_sched_gen_0_enable,
  input logic [15:0] strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides,
  input logic strg_ub_agg_only_agg_write_sched_gen_1_enable,
  input logic [15:0] strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides,
  input logic [3:0] strg_ub_agg_only_loops_in2buf_0_dimensionality,
  input logic [5:0] [15:0] strg_ub_agg_only_loops_in2buf_0_ranges,
  input logic [3:0] strg_ub_agg_only_loops_in2buf_1_dimensionality,
  input logic [5:0] [15:0] strg_ub_agg_only_loops_in2buf_1_ranges,
  input logic strg_ub_agg_sram_shared_agg_read_sched_gen_0_enable,
  input logic [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides,
  input logic strg_ub_agg_sram_shared_agg_read_sched_gen_1_enable,
  input logic [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides,
  input logic [3:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality,
  input logic [5:0] [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges,
  input logic [3:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality,
  input logic [5:0] [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges,
  input logic [8:0] strg_ub_sram_only_input_addr_gen_0_starting_addr,
  input logic [5:0] [8:0] strg_ub_sram_only_input_addr_gen_0_strides,
  input logic [8:0] strg_ub_sram_only_input_addr_gen_1_starting_addr,
  input logic [5:0] [8:0] strg_ub_sram_only_input_addr_gen_1_strides,
  input logic [8:0] strg_ub_sram_only_output_addr_gen_0_starting_addr,
  input logic [5:0] [8:0] strg_ub_sram_only_output_addr_gen_0_strides,
  input logic [8:0] strg_ub_sram_only_output_addr_gen_1_starting_addr,
  input logic [5:0] [8:0] strg_ub_sram_only_output_addr_gen_1_strides,
  input logic [3:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality,
  input logic [5:0] [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges,
  input logic [3:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality,
  input logic [5:0] [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges,
  input logic strg_ub_sram_tb_shared_output_sched_gen_0_enable,
  input logic [15:0] strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides,
  input logic strg_ub_sram_tb_shared_output_sched_gen_1_enable,
  input logic [15:0] strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides,
  input logic [3:0] strg_ub_tb_only_loops_buf2out_read_0_dimensionality,
  input logic [5:0] [15:0] strg_ub_tb_only_loops_buf2out_read_0_ranges,
  input logic [3:0] strg_ub_tb_only_loops_buf2out_read_1_dimensionality,
  input logic [5:0] [15:0] strg_ub_tb_only_loops_buf2out_read_1_ranges,
  input logic [3:0] strg_ub_tb_only_tb_read_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] strg_ub_tb_only_tb_read_addr_gen_0_strides,
  input logic [3:0] strg_ub_tb_only_tb_read_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] strg_ub_tb_only_tb_read_addr_gen_1_strides,
  input logic strg_ub_tb_only_tb_read_sched_gen_0_enable,
  input logic [15:0] strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides,
  input logic strg_ub_tb_only_tb_read_sched_gen_1_enable,
  input logic [15:0] strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides,
  input logic [3:0] strg_ub_tb_only_tb_write_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] strg_ub_tb_only_tb_write_addr_gen_0_strides,
  input logic [3:0] strg_ub_tb_only_tb_write_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] strg_ub_tb_only_tb_write_addr_gen_1_strides,
  input logic tile_en,
  input logic [1:0] wen_in,
  output logic [1:0] [31:0] config_data_out,
  output logic [1:0] [15:0] data_out,
  output logic empty,
  output logic full,
  output logic sram_ready_out,
  output logic stencil_valid,
  output logic [1:0] valid_out
);

logic [1:0] accessor_output;
logic [2:0][0:0][8:0] all_addr_to_mem;
logic [2:0][15:0] all_data_out;
logic [2:0][0:0][3:0][15:0] all_data_to_mem;
logic [2:0][0:0] all_ren_to_mem;
logic [2:0] all_valid_out;
logic [2:0][0:0] all_wen_to_mem;
logic cfg_seq_clk;
logic [1:0] chain_accessor_output;
logic [15:0] config_data_in_shrt;
logic [1:0][15:0] config_data_out_shrt;
logic config_seq_clk;
logic config_seq_clk_en;
logic [15:0] cycle_count;
logic [1:0][15:0] data_out_tile;
logic [0:0][8:0] fifo_addr_to_mem;
logic fifo_ctrl_clk;
logic [15:0] fifo_ctrl_data_in;
logic fifo_ctrl_pop;
logic fifo_ctrl_push;
logic [15:0] fifo_data_out;
logic [0:0][3:0][15:0] fifo_data_to_mem;
logic fifo_empty;
logic fifo_full;
logic fifo_ren_to_mem;
logic fifo_valid_out;
logic fifo_wen_to_mem;
logic gclk;
logic [2:0] loops_stencil_valid_mux_sel_out;
logic loops_stencil_valid_restart;
logic mem_0_clk;
logic mem_0_clk_en;
logic [8:0] mem_0_mem_addr_in_bank;
logic mem_0_mem_cen_in_bank;
logic [3:0][15:0] mem_0_mem_data_in_bank;
logic [0:0][3:0][15:0] mem_0_mem_data_out_bank;
logic mem_0_mem_wen_in_bank;
logic [8:0] mem_addr_cfg;
logic [0:0][0:0][8:0] mem_addr_dp;
logic [0:0][0:0][8:0] mem_addr_in;
logic [0:0] mem_cen_dp;
logic [0:0] mem_cen_in;
logic [3:0][15:0] mem_data_cfg;
logic [0:0][0:0][3:0][15:0] mem_data_dp;
logic [0:0][0:0][3:0][15:0] mem_data_in;
logic [0:0][3:0][15:0] mem_data_low_pt;
logic [0:0][0:0][3:0][15:0] mem_data_out;
logic mem_ren_cfg;
logic mem_wen_cfg;
logic [0:0] mem_wen_dp;
logic [0:0] mem_wen_in;
logic [1:0] mode_mask;
logic [0:0][8:0] sram_addr_to_mem;
logic sram_ctrl_clk;
logic [15:0] sram_ctrl_data_in;
logic [15:0] sram_ctrl_rd_addr_in;
logic sram_ctrl_ren;
logic sram_ctrl_wen;
logic [15:0] sram_ctrl_wr_addr_in;
logic [15:0] sram_data_out;
logic [0:0][3:0][15:0] sram_data_to_mem;
logic sram_ren_to_mem;
logic sram_valid_out;
logic sram_wen_to_mem;
logic stencil_valid_internal;
logic strg_ub_clk;
logic [0:0][0:0][8:0] ub_addr_to_mem;
logic [0:0] ub_cen_to_mem;
logic [1:0][15:0] ub_data_out;
logic [0:0][0:0][3:0][15:0] ub_data_to_mem;
logic [1:0] ub_valid_out;
logic [0:0] ub_wen_to_mem;
assign config_data_in_shrt = config_data_in[15:0];

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    cycle_count <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      cycle_count <= 16'h0;
    end
    else cycle_count <= cycle_count + 16'h1;
  end
end
assign stencil_valid = stencil_valid_internal;
assign config_data_out[0] = 32'(config_data_out_shrt[0]);
assign config_data_out[1] = 32'(config_data_out_shrt[1]);
assign gclk = clk & tile_en;
assign mem_data_low_pt[0] = mem_data_out[0][0];
assign cfg_seq_clk = gclk;
assign config_seq_clk = cfg_seq_clk;
assign config_seq_clk_en = clk_en | (|config_en);
assign mem_wen_in = (|config_en) ? mem_wen_cfg: mem_wen_dp;
assign mem_cen_in = (|config_en) ? mem_wen_cfg | mem_ren_cfg: mem_cen_dp;
assign mem_addr_in[0][0] = (|config_en) ? mem_addr_cfg: mem_addr_dp[0][0];
assign mem_data_in[0][0] = (|config_en) ? mem_data_cfg: mem_data_dp[0][0];
assign strg_ub_clk = gclk;
assign sram_ctrl_clk = gclk;
assign sram_ctrl_wen = wen_in[0];
assign sram_ctrl_ren = ren_in[0];
assign sram_ctrl_data_in = data_in[0];
assign sram_ctrl_wr_addr_in = addr_in[0];
assign sram_ctrl_rd_addr_in = addr_in[0];
assign fifo_ctrl_clk = gclk;
assign fifo_ctrl_data_in = data_in[0];
assign fifo_ctrl_push = wen_in[0];
assign fifo_ctrl_pop = ren_in[0];
assign empty = fifo_empty;
assign full = fifo_full;
assign all_data_to_mem[0] = ub_data_to_mem;
assign all_wen_to_mem[0] = ub_wen_to_mem;
assign all_ren_to_mem[0] = ub_cen_to_mem;
assign all_addr_to_mem[0] = ub_addr_to_mem;
assign all_data_to_mem[1] = fifo_data_to_mem;
assign all_wen_to_mem[1] = fifo_wen_to_mem;
assign all_ren_to_mem[1] = fifo_ren_to_mem;
assign all_addr_to_mem[1][0] = fifo_addr_to_mem[0];
assign all_data_to_mem[2] = sram_data_to_mem;
assign all_wen_to_mem[2] = sram_wen_to_mem;
assign all_ren_to_mem[2] = sram_ren_to_mem;
assign all_addr_to_mem[2][0] = sram_addr_to_mem[0];
assign mem_data_dp = all_data_to_mem[mode];
assign mem_cen_dp = all_ren_to_mem[mode] | all_wen_to_mem[mode];
assign mem_wen_dp = all_wen_to_mem[mode];
assign mem_addr_dp = all_addr_to_mem[mode];
assign mem_0_clk = gclk;
assign mem_0_clk_en = clk_en | (|config_en);
assign mem_0_mem_data_in_bank = mem_data_in[0];
assign mem_data_out[0] = mem_0_mem_data_out_bank;
assign mem_0_mem_addr_in_bank = mem_addr_in[0];
assign mem_0_mem_cen_in_bank = mem_cen_in;
assign mem_0_mem_wen_in_bank = mem_wen_in;
assign all_data_out[0] = ub_data_out[0];
assign all_valid_out[0] = ub_valid_out[0];
assign all_data_out[1] = fifo_data_out;
assign all_valid_out[1] = fifo_valid_out;
assign all_data_out[2] = sram_data_out;
assign all_valid_out[2] = sram_valid_out;
assign data_out_tile[0] = all_data_out[mode];
assign valid_out[0] = all_valid_out[mode];
assign data_out_tile[1] = ub_data_out[1];
assign valid_out[1] = ub_valid_out[1];
assign mode_mask[0] = |mode;
assign mode_mask[1] = 1'h0;
assign chain_accessor_output = accessor_output | mode_mask;
for_loop_6_16 #(
  .CONFIG_WIDTH(5'h10),
  .ITERATOR_SUPPORT(4'h6))
loops_stencil_valid (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_stencil_valid_dimensionality),
  .flush(flush),
  .ranges(loops_stencil_valid_ranges),
  .rst_n(rst_n),
  .step(stencil_valid_internal),
  .mux_sel_out(loops_stencil_valid_mux_sel_out),
  .restart(loops_stencil_valid_restart)
);

sched_gen_6_16 stencil_valid_sched_gen (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(stencil_valid_sched_gen_enable),
  .finished(loops_stencil_valid_restart),
  .flush(flush),
  .mux_sel(loops_stencil_valid_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(stencil_valid_sched_gen_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides(stencil_valid_sched_gen_sched_addr_gen_strides),
  .valid_output(stencil_valid_internal)
);

storage_config_seq config_seq (
  .clk(config_seq_clk),
  .clk_en(config_seq_clk_en),
  .config_addr_in(config_addr_in),
  .config_data_in(config_data_in_shrt),
  .config_en(config_en),
  .config_rd(config_read),
  .config_wr(config_write),
  .flush(flush),
  .rd_data_stg(mem_data_low_pt),
  .rst_n(rst_n),
  .addr_out(mem_addr_cfg),
  .rd_data_out(config_data_out_shrt),
  .ren_out(mem_ren_cfg),
  .wen_out(mem_wen_cfg),
  .wr_data(mem_data_cfg)
);

strg_ub_vec strg_ub (
  .agg_only_agg_read_addr_gen_0_starting_addr(strg_ub_agg_only_agg_read_addr_gen_0_starting_addr),
  .agg_only_agg_read_addr_gen_0_strides(strg_ub_agg_only_agg_read_addr_gen_0_strides),
  .agg_only_agg_read_addr_gen_1_starting_addr(strg_ub_agg_only_agg_read_addr_gen_1_starting_addr),
  .agg_only_agg_read_addr_gen_1_strides(strg_ub_agg_only_agg_read_addr_gen_1_strides),
  .agg_only_agg_write_addr_gen_0_starting_addr(strg_ub_agg_only_agg_write_addr_gen_0_starting_addr),
  .agg_only_agg_write_addr_gen_0_strides(strg_ub_agg_only_agg_write_addr_gen_0_strides),
  .agg_only_agg_write_addr_gen_1_starting_addr(strg_ub_agg_only_agg_write_addr_gen_1_starting_addr),
  .agg_only_agg_write_addr_gen_1_strides(strg_ub_agg_only_agg_write_addr_gen_1_strides),
  .agg_only_agg_write_sched_gen_0_enable(strg_ub_agg_only_agg_write_sched_gen_0_enable),
  .agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr),
  .agg_only_agg_write_sched_gen_0_sched_addr_gen_strides(strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides),
  .agg_only_agg_write_sched_gen_1_enable(strg_ub_agg_only_agg_write_sched_gen_1_enable),
  .agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr),
  .agg_only_agg_write_sched_gen_1_sched_addr_gen_strides(strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides),
  .agg_only_loops_in2buf_0_dimensionality(strg_ub_agg_only_loops_in2buf_0_dimensionality),
  .agg_only_loops_in2buf_0_ranges(strg_ub_agg_only_loops_in2buf_0_ranges),
  .agg_only_loops_in2buf_1_dimensionality(strg_ub_agg_only_loops_in2buf_1_dimensionality),
  .agg_only_loops_in2buf_1_ranges(strg_ub_agg_only_loops_in2buf_1_ranges),
  .agg_sram_shared_agg_read_sched_gen_0_enable(strg_ub_agg_sram_shared_agg_read_sched_gen_0_enable),
  .agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr),
  .agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides(strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides),
  .agg_sram_shared_agg_read_sched_gen_1_enable(strg_ub_agg_sram_shared_agg_read_sched_gen_1_enable),
  .agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr),
  .agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides(strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides),
  .agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality),
  .agg_sram_shared_loops_in2buf_autovec_write_0_ranges(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges),
  .agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality),
  .agg_sram_shared_loops_in2buf_autovec_write_1_ranges(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges),
  .clk(strg_ub_clk),
  .clk_en(clk_en),
  .data_from_strg(mem_data_out),
  .data_in(data_in),
  .flush(flush),
  .rst_n(rst_n),
  .sram_only_input_addr_gen_0_starting_addr(strg_ub_sram_only_input_addr_gen_0_starting_addr),
  .sram_only_input_addr_gen_0_strides(strg_ub_sram_only_input_addr_gen_0_strides),
  .sram_only_input_addr_gen_1_starting_addr(strg_ub_sram_only_input_addr_gen_1_starting_addr),
  .sram_only_input_addr_gen_1_strides(strg_ub_sram_only_input_addr_gen_1_strides),
  .sram_only_output_addr_gen_0_starting_addr(strg_ub_sram_only_output_addr_gen_0_starting_addr),
  .sram_only_output_addr_gen_0_strides(strg_ub_sram_only_output_addr_gen_0_strides),
  .sram_only_output_addr_gen_1_starting_addr(strg_ub_sram_only_output_addr_gen_1_starting_addr),
  .sram_only_output_addr_gen_1_strides(strg_ub_sram_only_output_addr_gen_1_strides),
  .sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality),
  .sram_tb_shared_loops_buf2out_autovec_read_0_ranges(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges),
  .sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality),
  .sram_tb_shared_loops_buf2out_autovec_read_1_ranges(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges),
  .sram_tb_shared_output_sched_gen_0_enable(strg_ub_sram_tb_shared_output_sched_gen_0_enable),
  .sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr),
  .sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides(strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides),
  .sram_tb_shared_output_sched_gen_1_enable(strg_ub_sram_tb_shared_output_sched_gen_1_enable),
  .sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr),
  .sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides(strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides),
  .tb_only_loops_buf2out_read_0_dimensionality(strg_ub_tb_only_loops_buf2out_read_0_dimensionality),
  .tb_only_loops_buf2out_read_0_ranges(strg_ub_tb_only_loops_buf2out_read_0_ranges),
  .tb_only_loops_buf2out_read_1_dimensionality(strg_ub_tb_only_loops_buf2out_read_1_dimensionality),
  .tb_only_loops_buf2out_read_1_ranges(strg_ub_tb_only_loops_buf2out_read_1_ranges),
  .tb_only_tb_read_addr_gen_0_starting_addr(strg_ub_tb_only_tb_read_addr_gen_0_starting_addr),
  .tb_only_tb_read_addr_gen_0_strides(strg_ub_tb_only_tb_read_addr_gen_0_strides),
  .tb_only_tb_read_addr_gen_1_starting_addr(strg_ub_tb_only_tb_read_addr_gen_1_starting_addr),
  .tb_only_tb_read_addr_gen_1_strides(strg_ub_tb_only_tb_read_addr_gen_1_strides),
  .tb_only_tb_read_sched_gen_0_enable(strg_ub_tb_only_tb_read_sched_gen_0_enable),
  .tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr),
  .tb_only_tb_read_sched_gen_0_sched_addr_gen_strides(strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides),
  .tb_only_tb_read_sched_gen_1_enable(strg_ub_tb_only_tb_read_sched_gen_1_enable),
  .tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr),
  .tb_only_tb_read_sched_gen_1_sched_addr_gen_strides(strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides),
  .tb_only_tb_write_addr_gen_0_starting_addr(strg_ub_tb_only_tb_write_addr_gen_0_starting_addr),
  .tb_only_tb_write_addr_gen_0_strides(strg_ub_tb_only_tb_write_addr_gen_0_strides),
  .tb_only_tb_write_addr_gen_1_starting_addr(strg_ub_tb_only_tb_write_addr_gen_1_starting_addr),
  .tb_only_tb_write_addr_gen_1_strides(strg_ub_tb_only_tb_write_addr_gen_1_strides),
  .accessor_output(accessor_output),
  .addr_out(ub_addr_to_mem),
  .cen_to_strg(ub_cen_to_mem),
  .data_out(ub_data_out),
  .data_to_strg(ub_data_to_mem),
  .wen_to_strg(ub_wen_to_mem)
);

strg_ram sram_ctrl (
  .clk(sram_ctrl_clk),
  .clk_en(clk_en),
  .data_from_strg(mem_data_out),
  .data_in(sram_ctrl_data_in),
  .flush(flush),
  .rd_addr_in(sram_ctrl_rd_addr_in),
  .ren(sram_ctrl_ren),
  .rst_n(rst_n),
  .wen(sram_ctrl_wen),
  .wr_addr_in(sram_ctrl_wr_addr_in),
  .addr_out(sram_addr_to_mem),
  .data_out(sram_data_out),
  .data_to_strg(sram_data_to_mem),
  .ready(sram_ready_out),
  .ren_to_strg(sram_ren_to_mem),
  .valid_out(sram_valid_out),
  .wen_to_strg(sram_wen_to_mem)
);

strg_fifo fifo_ctrl (
  .clk(fifo_ctrl_clk),
  .clk_en(clk_en),
  .data_from_strg(mem_data_out),
  .data_in(fifo_ctrl_data_in),
  .fifo_depth(fifo_ctrl_fifo_depth),
  .flush(flush),
  .pop(fifo_ctrl_pop),
  .push(fifo_ctrl_push),
  .rst_n(rst_n),
  .addr_out(fifo_addr_to_mem),
  .data_out(fifo_data_out),
  .data_to_strg(fifo_data_to_mem),
  .empty(fifo_empty),
  .full(fifo_full),
  .ren_to_strg(fifo_ren_to_mem),
  .valid_out(fifo_valid_out),
  .wen_to_strg(fifo_wen_to_mem)
);

TS1N16FFCLLSBLVTC512X32M4S_generator mem_0 (
  .clk(mem_0_clk),
  .clk_en(mem_0_clk_en),
  .flush(flush),
  .mem_addr_in_bank(mem_0_mem_addr_in_bank),
  .mem_cen_in_bank(mem_0_mem_cen_in_bank),
  .mem_data_in_bank(mem_0_mem_data_in_bank),
  .mem_wen_in_bank(mem_0_mem_wen_in_bank),
  .rtsel(2'h1),
  .wtsel(2'h0),
  .mem_data_out_bank(mem_0_mem_data_out_bank)
);

Chain chain (
  .accessor_output(chain_accessor_output),
  .chain_data_in(chain_data_in),
  .chain_en(chain_chain_en),
  .clk_en(clk_en),
  .curr_tile_data_out(data_out_tile),
  .flush(flush),
  .data_out_tile(data_out)
);

endmodule   // LakeTop

module LakeTop_W (
  input logic [15:0] addr_in_0,
  input logic [15:0] addr_in_1,
  input logic chain_chain_en,
  input logic [15:0] chain_data_in_0,
  input logic [15:0] chain_data_in_1,
  input logic clk,
  input logic clk_en,
  input logic [7:0] config_addr_in,
  input logic [31:0] config_data_in,
  input logic [1:0] config_en,
  input logic config_read,
  input logic config_write,
  input logic [15:0] data_in_0,
  input logic [15:0] data_in_1,
  input logic [15:0] fifo_ctrl_fifo_depth,
  input logic flush,
  input logic [3:0] loops_stencil_valid_dimensionality,
  input logic [15:0] loops_stencil_valid_ranges_0,
  input logic [15:0] loops_stencil_valid_ranges_1,
  input logic [15:0] loops_stencil_valid_ranges_2,
  input logic [15:0] loops_stencil_valid_ranges_3,
  input logic [15:0] loops_stencil_valid_ranges_4,
  input logic [15:0] loops_stencil_valid_ranges_5,
  input logic [1:0] mode,
  input logic [1:0] ren_in,
  input logic rst_n,
  input logic stencil_valid_sched_gen_enable,
  input logic [15:0] stencil_valid_sched_gen_sched_addr_gen_starting_addr,
  input logic [15:0] stencil_valid_sched_gen_sched_addr_gen_strides_0,
  input logic [15:0] stencil_valid_sched_gen_sched_addr_gen_strides_1,
  input logic [15:0] stencil_valid_sched_gen_sched_addr_gen_strides_2,
  input logic [15:0] stencil_valid_sched_gen_sched_addr_gen_strides_3,
  input logic [15:0] stencil_valid_sched_gen_sched_addr_gen_strides_4,
  input logic [15:0] stencil_valid_sched_gen_sched_addr_gen_strides_5,
  input logic [3:0] strg_ub_agg_only_agg_read_addr_gen_0_starting_addr,
  input logic [3:0] strg_ub_agg_only_agg_read_addr_gen_0_strides_0,
  input logic [3:0] strg_ub_agg_only_agg_read_addr_gen_0_strides_1,
  input logic [3:0] strg_ub_agg_only_agg_read_addr_gen_0_strides_2,
  input logic [3:0] strg_ub_agg_only_agg_read_addr_gen_0_strides_3,
  input logic [3:0] strg_ub_agg_only_agg_read_addr_gen_0_strides_4,
  input logic [3:0] strg_ub_agg_only_agg_read_addr_gen_0_strides_5,
  input logic [3:0] strg_ub_agg_only_agg_read_addr_gen_1_starting_addr,
  input logic [3:0] strg_ub_agg_only_agg_read_addr_gen_1_strides_0,
  input logic [3:0] strg_ub_agg_only_agg_read_addr_gen_1_strides_1,
  input logic [3:0] strg_ub_agg_only_agg_read_addr_gen_1_strides_2,
  input logic [3:0] strg_ub_agg_only_agg_read_addr_gen_1_strides_3,
  input logic [3:0] strg_ub_agg_only_agg_read_addr_gen_1_strides_4,
  input logic [3:0] strg_ub_agg_only_agg_read_addr_gen_1_strides_5,
  input logic [3:0] strg_ub_agg_only_agg_write_addr_gen_0_starting_addr,
  input logic [3:0] strg_ub_agg_only_agg_write_addr_gen_0_strides_0,
  input logic [3:0] strg_ub_agg_only_agg_write_addr_gen_0_strides_1,
  input logic [3:0] strg_ub_agg_only_agg_write_addr_gen_0_strides_2,
  input logic [3:0] strg_ub_agg_only_agg_write_addr_gen_0_strides_3,
  input logic [3:0] strg_ub_agg_only_agg_write_addr_gen_0_strides_4,
  input logic [3:0] strg_ub_agg_only_agg_write_addr_gen_0_strides_5,
  input logic [3:0] strg_ub_agg_only_agg_write_addr_gen_1_starting_addr,
  input logic [3:0] strg_ub_agg_only_agg_write_addr_gen_1_strides_0,
  input logic [3:0] strg_ub_agg_only_agg_write_addr_gen_1_strides_1,
  input logic [3:0] strg_ub_agg_only_agg_write_addr_gen_1_strides_2,
  input logic [3:0] strg_ub_agg_only_agg_write_addr_gen_1_strides_3,
  input logic [3:0] strg_ub_agg_only_agg_write_addr_gen_1_strides_4,
  input logic [3:0] strg_ub_agg_only_agg_write_addr_gen_1_strides_5,
  input logic strg_ub_agg_only_agg_write_sched_gen_0_enable,
  input logic [15:0] strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [15:0] strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0,
  input logic [15:0] strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1,
  input logic [15:0] strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2,
  input logic [15:0] strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3,
  input logic [15:0] strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4,
  input logic [15:0] strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5,
  input logic strg_ub_agg_only_agg_write_sched_gen_1_enable,
  input logic [15:0] strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [15:0] strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0,
  input logic [15:0] strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1,
  input logic [15:0] strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2,
  input logic [15:0] strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3,
  input logic [15:0] strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4,
  input logic [15:0] strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5,
  input logic [3:0] strg_ub_agg_only_loops_in2buf_0_dimensionality,
  input logic [15:0] strg_ub_agg_only_loops_in2buf_0_ranges_0,
  input logic [15:0] strg_ub_agg_only_loops_in2buf_0_ranges_1,
  input logic [15:0] strg_ub_agg_only_loops_in2buf_0_ranges_2,
  input logic [15:0] strg_ub_agg_only_loops_in2buf_0_ranges_3,
  input logic [15:0] strg_ub_agg_only_loops_in2buf_0_ranges_4,
  input logic [15:0] strg_ub_agg_only_loops_in2buf_0_ranges_5,
  input logic [3:0] strg_ub_agg_only_loops_in2buf_1_dimensionality,
  input logic [15:0] strg_ub_agg_only_loops_in2buf_1_ranges_0,
  input logic [15:0] strg_ub_agg_only_loops_in2buf_1_ranges_1,
  input logic [15:0] strg_ub_agg_only_loops_in2buf_1_ranges_2,
  input logic [15:0] strg_ub_agg_only_loops_in2buf_1_ranges_3,
  input logic [15:0] strg_ub_agg_only_loops_in2buf_1_ranges_4,
  input logic [15:0] strg_ub_agg_only_loops_in2buf_1_ranges_5,
  input logic strg_ub_agg_sram_shared_agg_read_sched_gen_0_enable,
  input logic [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0,
  input logic [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1,
  input logic [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2,
  input logic [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3,
  input logic [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4,
  input logic [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5,
  input logic strg_ub_agg_sram_shared_agg_read_sched_gen_1_enable,
  input logic [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0,
  input logic [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1,
  input logic [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2,
  input logic [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3,
  input logic [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4,
  input logic [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5,
  input logic [3:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality,
  input logic [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0,
  input logic [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1,
  input logic [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2,
  input logic [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3,
  input logic [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4,
  input logic [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5,
  input logic [3:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality,
  input logic [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0,
  input logic [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1,
  input logic [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2,
  input logic [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3,
  input logic [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4,
  input logic [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5,
  input logic [8:0] strg_ub_sram_only_input_addr_gen_0_starting_addr,
  input logic [8:0] strg_ub_sram_only_input_addr_gen_0_strides_0,
  input logic [8:0] strg_ub_sram_only_input_addr_gen_0_strides_1,
  input logic [8:0] strg_ub_sram_only_input_addr_gen_0_strides_2,
  input logic [8:0] strg_ub_sram_only_input_addr_gen_0_strides_3,
  input logic [8:0] strg_ub_sram_only_input_addr_gen_0_strides_4,
  input logic [8:0] strg_ub_sram_only_input_addr_gen_0_strides_5,
  input logic [8:0] strg_ub_sram_only_input_addr_gen_1_starting_addr,
  input logic [8:0] strg_ub_sram_only_input_addr_gen_1_strides_0,
  input logic [8:0] strg_ub_sram_only_input_addr_gen_1_strides_1,
  input logic [8:0] strg_ub_sram_only_input_addr_gen_1_strides_2,
  input logic [8:0] strg_ub_sram_only_input_addr_gen_1_strides_3,
  input logic [8:0] strg_ub_sram_only_input_addr_gen_1_strides_4,
  input logic [8:0] strg_ub_sram_only_input_addr_gen_1_strides_5,
  input logic [8:0] strg_ub_sram_only_output_addr_gen_0_starting_addr,
  input logic [8:0] strg_ub_sram_only_output_addr_gen_0_strides_0,
  input logic [8:0] strg_ub_sram_only_output_addr_gen_0_strides_1,
  input logic [8:0] strg_ub_sram_only_output_addr_gen_0_strides_2,
  input logic [8:0] strg_ub_sram_only_output_addr_gen_0_strides_3,
  input logic [8:0] strg_ub_sram_only_output_addr_gen_0_strides_4,
  input logic [8:0] strg_ub_sram_only_output_addr_gen_0_strides_5,
  input logic [8:0] strg_ub_sram_only_output_addr_gen_1_starting_addr,
  input logic [8:0] strg_ub_sram_only_output_addr_gen_1_strides_0,
  input logic [8:0] strg_ub_sram_only_output_addr_gen_1_strides_1,
  input logic [8:0] strg_ub_sram_only_output_addr_gen_1_strides_2,
  input logic [8:0] strg_ub_sram_only_output_addr_gen_1_strides_3,
  input logic [8:0] strg_ub_sram_only_output_addr_gen_1_strides_4,
  input logic [8:0] strg_ub_sram_only_output_addr_gen_1_strides_5,
  input logic [3:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality,
  input logic [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0,
  input logic [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1,
  input logic [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2,
  input logic [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3,
  input logic [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4,
  input logic [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5,
  input logic [3:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality,
  input logic [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0,
  input logic [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1,
  input logic [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2,
  input logic [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3,
  input logic [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4,
  input logic [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5,
  input logic strg_ub_sram_tb_shared_output_sched_gen_0_enable,
  input logic [15:0] strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [15:0] strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0,
  input logic [15:0] strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1,
  input logic [15:0] strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2,
  input logic [15:0] strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3,
  input logic [15:0] strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4,
  input logic [15:0] strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5,
  input logic strg_ub_sram_tb_shared_output_sched_gen_1_enable,
  input logic [15:0] strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [15:0] strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0,
  input logic [15:0] strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1,
  input logic [15:0] strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2,
  input logic [15:0] strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3,
  input logic [15:0] strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4,
  input logic [15:0] strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5,
  input logic [3:0] strg_ub_tb_only_loops_buf2out_read_0_dimensionality,
  input logic [15:0] strg_ub_tb_only_loops_buf2out_read_0_ranges_0,
  input logic [15:0] strg_ub_tb_only_loops_buf2out_read_0_ranges_1,
  input logic [15:0] strg_ub_tb_only_loops_buf2out_read_0_ranges_2,
  input logic [15:0] strg_ub_tb_only_loops_buf2out_read_0_ranges_3,
  input logic [15:0] strg_ub_tb_only_loops_buf2out_read_0_ranges_4,
  input logic [15:0] strg_ub_tb_only_loops_buf2out_read_0_ranges_5,
  input logic [3:0] strg_ub_tb_only_loops_buf2out_read_1_dimensionality,
  input logic [15:0] strg_ub_tb_only_loops_buf2out_read_1_ranges_0,
  input logic [15:0] strg_ub_tb_only_loops_buf2out_read_1_ranges_1,
  input logic [15:0] strg_ub_tb_only_loops_buf2out_read_1_ranges_2,
  input logic [15:0] strg_ub_tb_only_loops_buf2out_read_1_ranges_3,
  input logic [15:0] strg_ub_tb_only_loops_buf2out_read_1_ranges_4,
  input logic [15:0] strg_ub_tb_only_loops_buf2out_read_1_ranges_5,
  input logic [3:0] strg_ub_tb_only_tb_read_addr_gen_0_starting_addr,
  input logic [3:0] strg_ub_tb_only_tb_read_addr_gen_0_strides_0,
  input logic [3:0] strg_ub_tb_only_tb_read_addr_gen_0_strides_1,
  input logic [3:0] strg_ub_tb_only_tb_read_addr_gen_0_strides_2,
  input logic [3:0] strg_ub_tb_only_tb_read_addr_gen_0_strides_3,
  input logic [3:0] strg_ub_tb_only_tb_read_addr_gen_0_strides_4,
  input logic [3:0] strg_ub_tb_only_tb_read_addr_gen_0_strides_5,
  input logic [3:0] strg_ub_tb_only_tb_read_addr_gen_1_starting_addr,
  input logic [3:0] strg_ub_tb_only_tb_read_addr_gen_1_strides_0,
  input logic [3:0] strg_ub_tb_only_tb_read_addr_gen_1_strides_1,
  input logic [3:0] strg_ub_tb_only_tb_read_addr_gen_1_strides_2,
  input logic [3:0] strg_ub_tb_only_tb_read_addr_gen_1_strides_3,
  input logic [3:0] strg_ub_tb_only_tb_read_addr_gen_1_strides_4,
  input logic [3:0] strg_ub_tb_only_tb_read_addr_gen_1_strides_5,
  input logic strg_ub_tb_only_tb_read_sched_gen_0_enable,
  input logic [15:0] strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [15:0] strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0,
  input logic [15:0] strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1,
  input logic [15:0] strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2,
  input logic [15:0] strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3,
  input logic [15:0] strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4,
  input logic [15:0] strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5,
  input logic strg_ub_tb_only_tb_read_sched_gen_1_enable,
  input logic [15:0] strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [15:0] strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0,
  input logic [15:0] strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1,
  input logic [15:0] strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2,
  input logic [15:0] strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3,
  input logic [15:0] strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4,
  input logic [15:0] strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5,
  input logic [3:0] strg_ub_tb_only_tb_write_addr_gen_0_starting_addr,
  input logic [3:0] strg_ub_tb_only_tb_write_addr_gen_0_strides_0,
  input logic [3:0] strg_ub_tb_only_tb_write_addr_gen_0_strides_1,
  input logic [3:0] strg_ub_tb_only_tb_write_addr_gen_0_strides_2,
  input logic [3:0] strg_ub_tb_only_tb_write_addr_gen_0_strides_3,
  input logic [3:0] strg_ub_tb_only_tb_write_addr_gen_0_strides_4,
  input logic [3:0] strg_ub_tb_only_tb_write_addr_gen_0_strides_5,
  input logic [3:0] strg_ub_tb_only_tb_write_addr_gen_1_starting_addr,
  input logic [3:0] strg_ub_tb_only_tb_write_addr_gen_1_strides_0,
  input logic [3:0] strg_ub_tb_only_tb_write_addr_gen_1_strides_1,
  input logic [3:0] strg_ub_tb_only_tb_write_addr_gen_1_strides_2,
  input logic [3:0] strg_ub_tb_only_tb_write_addr_gen_1_strides_3,
  input logic [3:0] strg_ub_tb_only_tb_write_addr_gen_1_strides_4,
  input logic [3:0] strg_ub_tb_only_tb_write_addr_gen_1_strides_5,
  input logic tile_en,
  input logic [1:0] wen_in,
  output logic [31:0] config_data_out_0,
  output logic [31:0] config_data_out_1,
  output logic [15:0] data_out_0,
  output logic [15:0] data_out_1,
  output logic empty,
  output logic full,
  output logic sram_ready_out,
  output logic stencil_valid,
  output logic [1:0] valid_out
);

logic [1:0][15:0] LakeTop_addr_in;
logic [1:0][15:0] LakeTop_chain_data_in;
logic [1:0][31:0] LakeTop_config_data_out;
logic [1:0][15:0] LakeTop_data_in;
logic [1:0][15:0] LakeTop_data_out;
logic [5:0][15:0] LakeTop_loops_stencil_valid_ranges;
logic [5:0][15:0] LakeTop_stencil_valid_sched_gen_sched_addr_gen_strides;
logic [5:0][3:0] LakeTop_strg_ub_agg_only_agg_read_addr_gen_0_strides;
logic [5:0][3:0] LakeTop_strg_ub_agg_only_agg_read_addr_gen_1_strides;
logic [5:0][3:0] LakeTop_strg_ub_agg_only_agg_write_addr_gen_0_strides;
logic [5:0][3:0] LakeTop_strg_ub_agg_only_agg_write_addr_gen_1_strides;
logic [5:0][15:0] LakeTop_strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides;
logic [5:0][15:0] LakeTop_strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides;
logic [5:0][15:0] LakeTop_strg_ub_agg_only_loops_in2buf_0_ranges;
logic [5:0][15:0] LakeTop_strg_ub_agg_only_loops_in2buf_1_ranges;
logic [5:0][15:0] LakeTop_strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides;
logic [5:0][15:0] LakeTop_strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides;
logic [5:0][15:0] LakeTop_strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges;
logic [5:0][15:0] LakeTop_strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges;
logic [5:0][8:0] LakeTop_strg_ub_sram_only_input_addr_gen_0_strides;
logic [5:0][8:0] LakeTop_strg_ub_sram_only_input_addr_gen_1_strides;
logic [5:0][8:0] LakeTop_strg_ub_sram_only_output_addr_gen_0_strides;
logic [5:0][8:0] LakeTop_strg_ub_sram_only_output_addr_gen_1_strides;
logic [5:0][15:0] LakeTop_strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges;
logic [5:0][15:0] LakeTop_strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges;
logic [5:0][15:0] LakeTop_strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides;
logic [5:0][15:0] LakeTop_strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides;
logic [5:0][15:0] LakeTop_strg_ub_tb_only_loops_buf2out_read_0_ranges;
logic [5:0][15:0] LakeTop_strg_ub_tb_only_loops_buf2out_read_1_ranges;
logic [5:0][3:0] LakeTop_strg_ub_tb_only_tb_read_addr_gen_0_strides;
logic [5:0][3:0] LakeTop_strg_ub_tb_only_tb_read_addr_gen_1_strides;
logic [5:0][15:0] LakeTop_strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides;
logic [5:0][15:0] LakeTop_strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides;
logic [5:0][3:0] LakeTop_strg_ub_tb_only_tb_write_addr_gen_0_strides;
logic [5:0][3:0] LakeTop_strg_ub_tb_only_tb_write_addr_gen_1_strides;
assign LakeTop_addr_in[0] = addr_in_0;
assign LakeTop_addr_in[1] = addr_in_1;
assign LakeTop_chain_data_in[0] = chain_data_in_0;
assign LakeTop_chain_data_in[1] = chain_data_in_1;
assign config_data_out_0 = LakeTop_config_data_out[0];
assign config_data_out_1 = LakeTop_config_data_out[1];
assign LakeTop_data_in[0] = data_in_0;
assign LakeTop_data_in[1] = data_in_1;
assign data_out_0 = LakeTop_data_out[0];
assign data_out_1 = LakeTop_data_out[1];
assign LakeTop_loops_stencil_valid_ranges[0] = loops_stencil_valid_ranges_0;
assign LakeTop_loops_stencil_valid_ranges[1] = loops_stencil_valid_ranges_1;
assign LakeTop_loops_stencil_valid_ranges[2] = loops_stencil_valid_ranges_2;
assign LakeTop_loops_stencil_valid_ranges[3] = loops_stencil_valid_ranges_3;
assign LakeTop_loops_stencil_valid_ranges[4] = loops_stencil_valid_ranges_4;
assign LakeTop_loops_stencil_valid_ranges[5] = loops_stencil_valid_ranges_5;
assign LakeTop_stencil_valid_sched_gen_sched_addr_gen_strides[0] = stencil_valid_sched_gen_sched_addr_gen_strides_0;
assign LakeTop_stencil_valid_sched_gen_sched_addr_gen_strides[1] = stencil_valid_sched_gen_sched_addr_gen_strides_1;
assign LakeTop_stencil_valid_sched_gen_sched_addr_gen_strides[2] = stencil_valid_sched_gen_sched_addr_gen_strides_2;
assign LakeTop_stencil_valid_sched_gen_sched_addr_gen_strides[3] = stencil_valid_sched_gen_sched_addr_gen_strides_3;
assign LakeTop_stencil_valid_sched_gen_sched_addr_gen_strides[4] = stencil_valid_sched_gen_sched_addr_gen_strides_4;
assign LakeTop_stencil_valid_sched_gen_sched_addr_gen_strides[5] = stencil_valid_sched_gen_sched_addr_gen_strides_5;
assign LakeTop_strg_ub_agg_only_agg_read_addr_gen_0_strides[0] = strg_ub_agg_only_agg_read_addr_gen_0_strides_0;
assign LakeTop_strg_ub_agg_only_agg_read_addr_gen_0_strides[1] = strg_ub_agg_only_agg_read_addr_gen_0_strides_1;
assign LakeTop_strg_ub_agg_only_agg_read_addr_gen_0_strides[2] = strg_ub_agg_only_agg_read_addr_gen_0_strides_2;
assign LakeTop_strg_ub_agg_only_agg_read_addr_gen_0_strides[3] = strg_ub_agg_only_agg_read_addr_gen_0_strides_3;
assign LakeTop_strg_ub_agg_only_agg_read_addr_gen_0_strides[4] = strg_ub_agg_only_agg_read_addr_gen_0_strides_4;
assign LakeTop_strg_ub_agg_only_agg_read_addr_gen_0_strides[5] = strg_ub_agg_only_agg_read_addr_gen_0_strides_5;
assign LakeTop_strg_ub_agg_only_agg_read_addr_gen_1_strides[0] = strg_ub_agg_only_agg_read_addr_gen_1_strides_0;
assign LakeTop_strg_ub_agg_only_agg_read_addr_gen_1_strides[1] = strg_ub_agg_only_agg_read_addr_gen_1_strides_1;
assign LakeTop_strg_ub_agg_only_agg_read_addr_gen_1_strides[2] = strg_ub_agg_only_agg_read_addr_gen_1_strides_2;
assign LakeTop_strg_ub_agg_only_agg_read_addr_gen_1_strides[3] = strg_ub_agg_only_agg_read_addr_gen_1_strides_3;
assign LakeTop_strg_ub_agg_only_agg_read_addr_gen_1_strides[4] = strg_ub_agg_only_agg_read_addr_gen_1_strides_4;
assign LakeTop_strg_ub_agg_only_agg_read_addr_gen_1_strides[5] = strg_ub_agg_only_agg_read_addr_gen_1_strides_5;
assign LakeTop_strg_ub_agg_only_agg_write_addr_gen_0_strides[0] = strg_ub_agg_only_agg_write_addr_gen_0_strides_0;
assign LakeTop_strg_ub_agg_only_agg_write_addr_gen_0_strides[1] = strg_ub_agg_only_agg_write_addr_gen_0_strides_1;
assign LakeTop_strg_ub_agg_only_agg_write_addr_gen_0_strides[2] = strg_ub_agg_only_agg_write_addr_gen_0_strides_2;
assign LakeTop_strg_ub_agg_only_agg_write_addr_gen_0_strides[3] = strg_ub_agg_only_agg_write_addr_gen_0_strides_3;
assign LakeTop_strg_ub_agg_only_agg_write_addr_gen_0_strides[4] = strg_ub_agg_only_agg_write_addr_gen_0_strides_4;
assign LakeTop_strg_ub_agg_only_agg_write_addr_gen_0_strides[5] = strg_ub_agg_only_agg_write_addr_gen_0_strides_5;
assign LakeTop_strg_ub_agg_only_agg_write_addr_gen_1_strides[0] = strg_ub_agg_only_agg_write_addr_gen_1_strides_0;
assign LakeTop_strg_ub_agg_only_agg_write_addr_gen_1_strides[1] = strg_ub_agg_only_agg_write_addr_gen_1_strides_1;
assign LakeTop_strg_ub_agg_only_agg_write_addr_gen_1_strides[2] = strg_ub_agg_only_agg_write_addr_gen_1_strides_2;
assign LakeTop_strg_ub_agg_only_agg_write_addr_gen_1_strides[3] = strg_ub_agg_only_agg_write_addr_gen_1_strides_3;
assign LakeTop_strg_ub_agg_only_agg_write_addr_gen_1_strides[4] = strg_ub_agg_only_agg_write_addr_gen_1_strides_4;
assign LakeTop_strg_ub_agg_only_agg_write_addr_gen_1_strides[5] = strg_ub_agg_only_agg_write_addr_gen_1_strides_5;
assign LakeTop_strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides[0] = strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0;
assign LakeTop_strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides[1] = strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1;
assign LakeTop_strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides[2] = strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2;
assign LakeTop_strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides[3] = strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3;
assign LakeTop_strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides[4] = strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4;
assign LakeTop_strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides[5] = strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5;
assign LakeTop_strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides[0] = strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0;
assign LakeTop_strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides[1] = strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1;
assign LakeTop_strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides[2] = strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2;
assign LakeTop_strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides[3] = strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3;
assign LakeTop_strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides[4] = strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4;
assign LakeTop_strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides[5] = strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5;
assign LakeTop_strg_ub_agg_only_loops_in2buf_0_ranges[0] = strg_ub_agg_only_loops_in2buf_0_ranges_0;
assign LakeTop_strg_ub_agg_only_loops_in2buf_0_ranges[1] = strg_ub_agg_only_loops_in2buf_0_ranges_1;
assign LakeTop_strg_ub_agg_only_loops_in2buf_0_ranges[2] = strg_ub_agg_only_loops_in2buf_0_ranges_2;
assign LakeTop_strg_ub_agg_only_loops_in2buf_0_ranges[3] = strg_ub_agg_only_loops_in2buf_0_ranges_3;
assign LakeTop_strg_ub_agg_only_loops_in2buf_0_ranges[4] = strg_ub_agg_only_loops_in2buf_0_ranges_4;
assign LakeTop_strg_ub_agg_only_loops_in2buf_0_ranges[5] = strg_ub_agg_only_loops_in2buf_0_ranges_5;
assign LakeTop_strg_ub_agg_only_loops_in2buf_1_ranges[0] = strg_ub_agg_only_loops_in2buf_1_ranges_0;
assign LakeTop_strg_ub_agg_only_loops_in2buf_1_ranges[1] = strg_ub_agg_only_loops_in2buf_1_ranges_1;
assign LakeTop_strg_ub_agg_only_loops_in2buf_1_ranges[2] = strg_ub_agg_only_loops_in2buf_1_ranges_2;
assign LakeTop_strg_ub_agg_only_loops_in2buf_1_ranges[3] = strg_ub_agg_only_loops_in2buf_1_ranges_3;
assign LakeTop_strg_ub_agg_only_loops_in2buf_1_ranges[4] = strg_ub_agg_only_loops_in2buf_1_ranges_4;
assign LakeTop_strg_ub_agg_only_loops_in2buf_1_ranges[5] = strg_ub_agg_only_loops_in2buf_1_ranges_5;
assign LakeTop_strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides[0] = strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0;
assign LakeTop_strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides[1] = strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1;
assign LakeTop_strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides[2] = strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2;
assign LakeTop_strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides[3] = strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3;
assign LakeTop_strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides[4] = strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4;
assign LakeTop_strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides[5] = strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5;
assign LakeTop_strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides[0] = strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0;
assign LakeTop_strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides[1] = strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1;
assign LakeTop_strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides[2] = strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2;
assign LakeTop_strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides[3] = strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3;
assign LakeTop_strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides[4] = strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4;
assign LakeTop_strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides[5] = strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5;
assign LakeTop_strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges[0] = strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0;
assign LakeTop_strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges[1] = strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1;
assign LakeTop_strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges[2] = strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2;
assign LakeTop_strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges[3] = strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3;
assign LakeTop_strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges[4] = strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4;
assign LakeTop_strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges[5] = strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5;
assign LakeTop_strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges[0] = strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0;
assign LakeTop_strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges[1] = strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1;
assign LakeTop_strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges[2] = strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2;
assign LakeTop_strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges[3] = strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3;
assign LakeTop_strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges[4] = strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4;
assign LakeTop_strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges[5] = strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5;
assign LakeTop_strg_ub_sram_only_input_addr_gen_0_strides[0] = strg_ub_sram_only_input_addr_gen_0_strides_0;
assign LakeTop_strg_ub_sram_only_input_addr_gen_0_strides[1] = strg_ub_sram_only_input_addr_gen_0_strides_1;
assign LakeTop_strg_ub_sram_only_input_addr_gen_0_strides[2] = strg_ub_sram_only_input_addr_gen_0_strides_2;
assign LakeTop_strg_ub_sram_only_input_addr_gen_0_strides[3] = strg_ub_sram_only_input_addr_gen_0_strides_3;
assign LakeTop_strg_ub_sram_only_input_addr_gen_0_strides[4] = strg_ub_sram_only_input_addr_gen_0_strides_4;
assign LakeTop_strg_ub_sram_only_input_addr_gen_0_strides[5] = strg_ub_sram_only_input_addr_gen_0_strides_5;
assign LakeTop_strg_ub_sram_only_input_addr_gen_1_strides[0] = strg_ub_sram_only_input_addr_gen_1_strides_0;
assign LakeTop_strg_ub_sram_only_input_addr_gen_1_strides[1] = strg_ub_sram_only_input_addr_gen_1_strides_1;
assign LakeTop_strg_ub_sram_only_input_addr_gen_1_strides[2] = strg_ub_sram_only_input_addr_gen_1_strides_2;
assign LakeTop_strg_ub_sram_only_input_addr_gen_1_strides[3] = strg_ub_sram_only_input_addr_gen_1_strides_3;
assign LakeTop_strg_ub_sram_only_input_addr_gen_1_strides[4] = strg_ub_sram_only_input_addr_gen_1_strides_4;
assign LakeTop_strg_ub_sram_only_input_addr_gen_1_strides[5] = strg_ub_sram_only_input_addr_gen_1_strides_5;
assign LakeTop_strg_ub_sram_only_output_addr_gen_0_strides[0] = strg_ub_sram_only_output_addr_gen_0_strides_0;
assign LakeTop_strg_ub_sram_only_output_addr_gen_0_strides[1] = strg_ub_sram_only_output_addr_gen_0_strides_1;
assign LakeTop_strg_ub_sram_only_output_addr_gen_0_strides[2] = strg_ub_sram_only_output_addr_gen_0_strides_2;
assign LakeTop_strg_ub_sram_only_output_addr_gen_0_strides[3] = strg_ub_sram_only_output_addr_gen_0_strides_3;
assign LakeTop_strg_ub_sram_only_output_addr_gen_0_strides[4] = strg_ub_sram_only_output_addr_gen_0_strides_4;
assign LakeTop_strg_ub_sram_only_output_addr_gen_0_strides[5] = strg_ub_sram_only_output_addr_gen_0_strides_5;
assign LakeTop_strg_ub_sram_only_output_addr_gen_1_strides[0] = strg_ub_sram_only_output_addr_gen_1_strides_0;
assign LakeTop_strg_ub_sram_only_output_addr_gen_1_strides[1] = strg_ub_sram_only_output_addr_gen_1_strides_1;
assign LakeTop_strg_ub_sram_only_output_addr_gen_1_strides[2] = strg_ub_sram_only_output_addr_gen_1_strides_2;
assign LakeTop_strg_ub_sram_only_output_addr_gen_1_strides[3] = strg_ub_sram_only_output_addr_gen_1_strides_3;
assign LakeTop_strg_ub_sram_only_output_addr_gen_1_strides[4] = strg_ub_sram_only_output_addr_gen_1_strides_4;
assign LakeTop_strg_ub_sram_only_output_addr_gen_1_strides[5] = strg_ub_sram_only_output_addr_gen_1_strides_5;
assign LakeTop_strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges[0] = strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0;
assign LakeTop_strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges[1] = strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1;
assign LakeTop_strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges[2] = strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2;
assign LakeTop_strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges[3] = strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3;
assign LakeTop_strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges[4] = strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4;
assign LakeTop_strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges[5] = strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5;
assign LakeTop_strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges[0] = strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0;
assign LakeTop_strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges[1] = strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1;
assign LakeTop_strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges[2] = strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2;
assign LakeTop_strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges[3] = strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3;
assign LakeTop_strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges[4] = strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4;
assign LakeTop_strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges[5] = strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5;
assign LakeTop_strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides[0] = strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0;
assign LakeTop_strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides[1] = strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1;
assign LakeTop_strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides[2] = strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2;
assign LakeTop_strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides[3] = strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3;
assign LakeTop_strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides[4] = strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4;
assign LakeTop_strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides[5] = strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5;
assign LakeTop_strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides[0] = strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0;
assign LakeTop_strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides[1] = strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1;
assign LakeTop_strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides[2] = strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2;
assign LakeTop_strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides[3] = strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3;
assign LakeTop_strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides[4] = strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4;
assign LakeTop_strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides[5] = strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5;
assign LakeTop_strg_ub_tb_only_loops_buf2out_read_0_ranges[0] = strg_ub_tb_only_loops_buf2out_read_0_ranges_0;
assign LakeTop_strg_ub_tb_only_loops_buf2out_read_0_ranges[1] = strg_ub_tb_only_loops_buf2out_read_0_ranges_1;
assign LakeTop_strg_ub_tb_only_loops_buf2out_read_0_ranges[2] = strg_ub_tb_only_loops_buf2out_read_0_ranges_2;
assign LakeTop_strg_ub_tb_only_loops_buf2out_read_0_ranges[3] = strg_ub_tb_only_loops_buf2out_read_0_ranges_3;
assign LakeTop_strg_ub_tb_only_loops_buf2out_read_0_ranges[4] = strg_ub_tb_only_loops_buf2out_read_0_ranges_4;
assign LakeTop_strg_ub_tb_only_loops_buf2out_read_0_ranges[5] = strg_ub_tb_only_loops_buf2out_read_0_ranges_5;
assign LakeTop_strg_ub_tb_only_loops_buf2out_read_1_ranges[0] = strg_ub_tb_only_loops_buf2out_read_1_ranges_0;
assign LakeTop_strg_ub_tb_only_loops_buf2out_read_1_ranges[1] = strg_ub_tb_only_loops_buf2out_read_1_ranges_1;
assign LakeTop_strg_ub_tb_only_loops_buf2out_read_1_ranges[2] = strg_ub_tb_only_loops_buf2out_read_1_ranges_2;
assign LakeTop_strg_ub_tb_only_loops_buf2out_read_1_ranges[3] = strg_ub_tb_only_loops_buf2out_read_1_ranges_3;
assign LakeTop_strg_ub_tb_only_loops_buf2out_read_1_ranges[4] = strg_ub_tb_only_loops_buf2out_read_1_ranges_4;
assign LakeTop_strg_ub_tb_only_loops_buf2out_read_1_ranges[5] = strg_ub_tb_only_loops_buf2out_read_1_ranges_5;
assign LakeTop_strg_ub_tb_only_tb_read_addr_gen_0_strides[0] = strg_ub_tb_only_tb_read_addr_gen_0_strides_0;
assign LakeTop_strg_ub_tb_only_tb_read_addr_gen_0_strides[1] = strg_ub_tb_only_tb_read_addr_gen_0_strides_1;
assign LakeTop_strg_ub_tb_only_tb_read_addr_gen_0_strides[2] = strg_ub_tb_only_tb_read_addr_gen_0_strides_2;
assign LakeTop_strg_ub_tb_only_tb_read_addr_gen_0_strides[3] = strg_ub_tb_only_tb_read_addr_gen_0_strides_3;
assign LakeTop_strg_ub_tb_only_tb_read_addr_gen_0_strides[4] = strg_ub_tb_only_tb_read_addr_gen_0_strides_4;
assign LakeTop_strg_ub_tb_only_tb_read_addr_gen_0_strides[5] = strg_ub_tb_only_tb_read_addr_gen_0_strides_5;
assign LakeTop_strg_ub_tb_only_tb_read_addr_gen_1_strides[0] = strg_ub_tb_only_tb_read_addr_gen_1_strides_0;
assign LakeTop_strg_ub_tb_only_tb_read_addr_gen_1_strides[1] = strg_ub_tb_only_tb_read_addr_gen_1_strides_1;
assign LakeTop_strg_ub_tb_only_tb_read_addr_gen_1_strides[2] = strg_ub_tb_only_tb_read_addr_gen_1_strides_2;
assign LakeTop_strg_ub_tb_only_tb_read_addr_gen_1_strides[3] = strg_ub_tb_only_tb_read_addr_gen_1_strides_3;
assign LakeTop_strg_ub_tb_only_tb_read_addr_gen_1_strides[4] = strg_ub_tb_only_tb_read_addr_gen_1_strides_4;
assign LakeTop_strg_ub_tb_only_tb_read_addr_gen_1_strides[5] = strg_ub_tb_only_tb_read_addr_gen_1_strides_5;
assign LakeTop_strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides[0] = strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0;
assign LakeTop_strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides[1] = strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1;
assign LakeTop_strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides[2] = strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2;
assign LakeTop_strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides[3] = strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3;
assign LakeTop_strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides[4] = strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4;
assign LakeTop_strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides[5] = strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5;
assign LakeTop_strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides[0] = strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0;
assign LakeTop_strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides[1] = strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1;
assign LakeTop_strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides[2] = strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2;
assign LakeTop_strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides[3] = strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3;
assign LakeTop_strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides[4] = strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4;
assign LakeTop_strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides[5] = strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5;
assign LakeTop_strg_ub_tb_only_tb_write_addr_gen_0_strides[0] = strg_ub_tb_only_tb_write_addr_gen_0_strides_0;
assign LakeTop_strg_ub_tb_only_tb_write_addr_gen_0_strides[1] = strg_ub_tb_only_tb_write_addr_gen_0_strides_1;
assign LakeTop_strg_ub_tb_only_tb_write_addr_gen_0_strides[2] = strg_ub_tb_only_tb_write_addr_gen_0_strides_2;
assign LakeTop_strg_ub_tb_only_tb_write_addr_gen_0_strides[3] = strg_ub_tb_only_tb_write_addr_gen_0_strides_3;
assign LakeTop_strg_ub_tb_only_tb_write_addr_gen_0_strides[4] = strg_ub_tb_only_tb_write_addr_gen_0_strides_4;
assign LakeTop_strg_ub_tb_only_tb_write_addr_gen_0_strides[5] = strg_ub_tb_only_tb_write_addr_gen_0_strides_5;
assign LakeTop_strg_ub_tb_only_tb_write_addr_gen_1_strides[0] = strg_ub_tb_only_tb_write_addr_gen_1_strides_0;
assign LakeTop_strg_ub_tb_only_tb_write_addr_gen_1_strides[1] = strg_ub_tb_only_tb_write_addr_gen_1_strides_1;
assign LakeTop_strg_ub_tb_only_tb_write_addr_gen_1_strides[2] = strg_ub_tb_only_tb_write_addr_gen_1_strides_2;
assign LakeTop_strg_ub_tb_only_tb_write_addr_gen_1_strides[3] = strg_ub_tb_only_tb_write_addr_gen_1_strides_3;
assign LakeTop_strg_ub_tb_only_tb_write_addr_gen_1_strides[4] = strg_ub_tb_only_tb_write_addr_gen_1_strides_4;
assign LakeTop_strg_ub_tb_only_tb_write_addr_gen_1_strides[5] = strg_ub_tb_only_tb_write_addr_gen_1_strides_5;
LakeTop LakeTop (
  .addr_in(LakeTop_addr_in),
  .chain_chain_en(chain_chain_en),
  .chain_data_in(LakeTop_chain_data_in),
  .clk(clk),
  .clk_en(clk_en),
  .config_addr_in(config_addr_in),
  .config_data_in(config_data_in),
  .config_en(config_en),
  .config_read(config_read),
  .config_write(config_write),
  .data_in(LakeTop_data_in),
  .fifo_ctrl_fifo_depth(fifo_ctrl_fifo_depth),
  .flush(flush),
  .loops_stencil_valid_dimensionality(loops_stencil_valid_dimensionality),
  .loops_stencil_valid_ranges(LakeTop_loops_stencil_valid_ranges),
  .mode(mode),
  .ren_in(ren_in),
  .rst_n(rst_n),
  .stencil_valid_sched_gen_enable(stencil_valid_sched_gen_enable),
  .stencil_valid_sched_gen_sched_addr_gen_starting_addr(stencil_valid_sched_gen_sched_addr_gen_starting_addr),
  .stencil_valid_sched_gen_sched_addr_gen_strides(LakeTop_stencil_valid_sched_gen_sched_addr_gen_strides),
  .strg_ub_agg_only_agg_read_addr_gen_0_starting_addr(strg_ub_agg_only_agg_read_addr_gen_0_starting_addr),
  .strg_ub_agg_only_agg_read_addr_gen_0_strides(LakeTop_strg_ub_agg_only_agg_read_addr_gen_0_strides),
  .strg_ub_agg_only_agg_read_addr_gen_1_starting_addr(strg_ub_agg_only_agg_read_addr_gen_1_starting_addr),
  .strg_ub_agg_only_agg_read_addr_gen_1_strides(LakeTop_strg_ub_agg_only_agg_read_addr_gen_1_strides),
  .strg_ub_agg_only_agg_write_addr_gen_0_starting_addr(strg_ub_agg_only_agg_write_addr_gen_0_starting_addr),
  .strg_ub_agg_only_agg_write_addr_gen_0_strides(LakeTop_strg_ub_agg_only_agg_write_addr_gen_0_strides),
  .strg_ub_agg_only_agg_write_addr_gen_1_starting_addr(strg_ub_agg_only_agg_write_addr_gen_1_starting_addr),
  .strg_ub_agg_only_agg_write_addr_gen_1_strides(LakeTop_strg_ub_agg_only_agg_write_addr_gen_1_strides),
  .strg_ub_agg_only_agg_write_sched_gen_0_enable(strg_ub_agg_only_agg_write_sched_gen_0_enable),
  .strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr),
  .strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides(LakeTop_strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides),
  .strg_ub_agg_only_agg_write_sched_gen_1_enable(strg_ub_agg_only_agg_write_sched_gen_1_enable),
  .strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr),
  .strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides(LakeTop_strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides),
  .strg_ub_agg_only_loops_in2buf_0_dimensionality(strg_ub_agg_only_loops_in2buf_0_dimensionality),
  .strg_ub_agg_only_loops_in2buf_0_ranges(LakeTop_strg_ub_agg_only_loops_in2buf_0_ranges),
  .strg_ub_agg_only_loops_in2buf_1_dimensionality(strg_ub_agg_only_loops_in2buf_1_dimensionality),
  .strg_ub_agg_only_loops_in2buf_1_ranges(LakeTop_strg_ub_agg_only_loops_in2buf_1_ranges),
  .strg_ub_agg_sram_shared_agg_read_sched_gen_0_enable(strg_ub_agg_sram_shared_agg_read_sched_gen_0_enable),
  .strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr),
  .strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides(LakeTop_strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides),
  .strg_ub_agg_sram_shared_agg_read_sched_gen_1_enable(strg_ub_agg_sram_shared_agg_read_sched_gen_1_enable),
  .strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr),
  .strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides(LakeTop_strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides),
  .strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality),
  .strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges(LakeTop_strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges),
  .strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality),
  .strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges(LakeTop_strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges),
  .strg_ub_sram_only_input_addr_gen_0_starting_addr(strg_ub_sram_only_input_addr_gen_0_starting_addr),
  .strg_ub_sram_only_input_addr_gen_0_strides(LakeTop_strg_ub_sram_only_input_addr_gen_0_strides),
  .strg_ub_sram_only_input_addr_gen_1_starting_addr(strg_ub_sram_only_input_addr_gen_1_starting_addr),
  .strg_ub_sram_only_input_addr_gen_1_strides(LakeTop_strg_ub_sram_only_input_addr_gen_1_strides),
  .strg_ub_sram_only_output_addr_gen_0_starting_addr(strg_ub_sram_only_output_addr_gen_0_starting_addr),
  .strg_ub_sram_only_output_addr_gen_0_strides(LakeTop_strg_ub_sram_only_output_addr_gen_0_strides),
  .strg_ub_sram_only_output_addr_gen_1_starting_addr(strg_ub_sram_only_output_addr_gen_1_starting_addr),
  .strg_ub_sram_only_output_addr_gen_1_strides(LakeTop_strg_ub_sram_only_output_addr_gen_1_strides),
  .strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality),
  .strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges(LakeTop_strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges),
  .strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality),
  .strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges(LakeTop_strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges),
  .strg_ub_sram_tb_shared_output_sched_gen_0_enable(strg_ub_sram_tb_shared_output_sched_gen_0_enable),
  .strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr),
  .strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides(LakeTop_strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides),
  .strg_ub_sram_tb_shared_output_sched_gen_1_enable(strg_ub_sram_tb_shared_output_sched_gen_1_enable),
  .strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr),
  .strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides(LakeTop_strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides),
  .strg_ub_tb_only_loops_buf2out_read_0_dimensionality(strg_ub_tb_only_loops_buf2out_read_0_dimensionality),
  .strg_ub_tb_only_loops_buf2out_read_0_ranges(LakeTop_strg_ub_tb_only_loops_buf2out_read_0_ranges),
  .strg_ub_tb_only_loops_buf2out_read_1_dimensionality(strg_ub_tb_only_loops_buf2out_read_1_dimensionality),
  .strg_ub_tb_only_loops_buf2out_read_1_ranges(LakeTop_strg_ub_tb_only_loops_buf2out_read_1_ranges),
  .strg_ub_tb_only_tb_read_addr_gen_0_starting_addr(strg_ub_tb_only_tb_read_addr_gen_0_starting_addr),
  .strg_ub_tb_only_tb_read_addr_gen_0_strides(LakeTop_strg_ub_tb_only_tb_read_addr_gen_0_strides),
  .strg_ub_tb_only_tb_read_addr_gen_1_starting_addr(strg_ub_tb_only_tb_read_addr_gen_1_starting_addr),
  .strg_ub_tb_only_tb_read_addr_gen_1_strides(LakeTop_strg_ub_tb_only_tb_read_addr_gen_1_strides),
  .strg_ub_tb_only_tb_read_sched_gen_0_enable(strg_ub_tb_only_tb_read_sched_gen_0_enable),
  .strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr),
  .strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides(LakeTop_strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides),
  .strg_ub_tb_only_tb_read_sched_gen_1_enable(strg_ub_tb_only_tb_read_sched_gen_1_enable),
  .strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr),
  .strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides(LakeTop_strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides),
  .strg_ub_tb_only_tb_write_addr_gen_0_starting_addr(strg_ub_tb_only_tb_write_addr_gen_0_starting_addr),
  .strg_ub_tb_only_tb_write_addr_gen_0_strides(LakeTop_strg_ub_tb_only_tb_write_addr_gen_0_strides),
  .strg_ub_tb_only_tb_write_addr_gen_1_starting_addr(strg_ub_tb_only_tb_write_addr_gen_1_starting_addr),
  .strg_ub_tb_only_tb_write_addr_gen_1_strides(LakeTop_strg_ub_tb_only_tb_write_addr_gen_1_strides),
  .tile_en(tile_en),
  .wen_in(wen_in),
  .config_data_out(LakeTop_config_data_out),
  .data_out(LakeTop_data_out),
  .empty(empty),
  .full(full),
  .sram_ready_out(sram_ready_out),
  .stencil_valid(stencil_valid),
  .valid_out(valid_out)
);

endmodule   // LakeTop_W

module TS1N16FFCLLSBLVTC512X32M4S_generator (
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [8:0] mem_addr_in_bank,
  input logic mem_cen_in_bank,
  input logic [3:0] [15:0] mem_data_in_bank,
  input logic mem_wen_in_bank,
  input logic [1:0] rtsel,
  input logic [1:0] wtsel,
  output logic [0:0][3:0] [15:0] mem_data_out_bank
);

logic [8:0] mem_addr_to_sram;
always_comb begin
  mem_addr_to_sram = mem_addr_in_bank;
end
sram_stub mem_0 (
  .addr(mem_addr_to_sram),
  .cen(mem_cen_in_bank),
  .clk(clk),
  .clk_en(clk_en),
  .data_in(mem_data_in_bank),
  .flush(flush),
  .wen(mem_wen_in_bank),
  .data_out(mem_data_out_bank)
);

endmodule   // TS1N16FFCLLSBLVTC512X32M4S_generator

module addr_gen_6_16 (
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [2:0] mux_sel,
  input logic restart,
  input logic rst_n,
  input logic [15:0] starting_addr,
  input logic step,
  input logic [5:0] [15:0] strides,
  output logic [15:0] addr_out
);

logic [15:0] calc_addr;
logic [15:0] current_addr;
logic [15:0] strt_addr;
assign strt_addr = starting_addr;
assign addr_out = calc_addr;
assign calc_addr = strt_addr + current_addr;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    current_addr <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      current_addr <= 16'h0;
    end
    else if (step) begin
      if (restart) begin
        current_addr <= 16'h0;
      end
      else current_addr <= current_addr + strides[mux_sel];
    end
  end
end
endmodule   // addr_gen_6_16

module addr_gen_6_4 (
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [2:0] mux_sel,
  input logic restart,
  input logic rst_n,
  input logic [3:0] starting_addr,
  input logic step,
  input logic [5:0] [3:0] strides,
  output logic [3:0] addr_out
);

logic [3:0] calc_addr;
logic [3:0] current_addr;
logic [3:0] strt_addr;
assign strt_addr = starting_addr;
assign addr_out = calc_addr;
assign calc_addr = strt_addr + current_addr;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    current_addr <= 4'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      current_addr <= 4'h0;
    end
    else if (step) begin
      if (restart) begin
        current_addr <= 4'h0;
      end
      else current_addr <= current_addr + strides[mux_sel];
    end
  end
end
endmodule   // addr_gen_6_4

module addr_gen_6_9 (
  input logic clk,
  input logic clk_en,
  input logic flush,
  input logic [2:0] mux_sel,
  input logic restart,
  input logic rst_n,
  input logic [8:0] starting_addr,
  input logic step,
  input logic [5:0] [8:0] strides,
  output logic [8:0] addr_out
);

logic [8:0] calc_addr;
logic [8:0] current_addr;
logic [8:0] strt_addr;
assign strt_addr = starting_addr;
assign addr_out = calc_addr;
assign calc_addr = strt_addr + current_addr;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    current_addr <= 9'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      current_addr <= 9'h0;
    end
    else if (step) begin
      if (restart) begin
        current_addr <= 9'h0;
      end
      else current_addr <= current_addr + strides[mux_sel];
    end
  end
end
endmodule   // addr_gen_6_9

module for_loop_6_16 #(
  parameter CONFIG_WIDTH = 5'h10,
  parameter ITERATOR_SUPPORT = 4'h6
)
(
  input logic clk,
  input logic clk_en,
  input logic [3:0] dimensionality,
  input logic flush,
  input logic [5:0] [15:0] ranges,
  input logic rst_n,
  input logic step,
  output logic [2:0] mux_sel_out,
  output logic restart
);

logic [5:0] clear;
logic [5:0][15:0] dim_counter;
logic done;
logic [5:0] inc;
logic [15:0] inced_cnt;
logic [5:0] max_value;
logic maxed_value;
logic [2:0] mux_sel;
assign mux_sel_out = mux_sel;
assign inced_cnt = dim_counter[mux_sel] + 16'h1;
assign maxed_value = (dim_counter[mux_sel] == ranges[mux_sel]) & inc[mux_sel];
always_comb begin
  mux_sel = 3'h0;
  done = 1'h0;
  if (~done) begin
    if ((~max_value[0]) & (dimensionality > 4'h0)) begin
      mux_sel = 3'h0;
      done = 1'h1;
    end
  end
  if (~done) begin
    if ((~max_value[1]) & (dimensionality > 4'h1)) begin
      mux_sel = 3'h1;
      done = 1'h1;
    end
  end
  if (~done) begin
    if ((~max_value[2]) & (dimensionality > 4'h2)) begin
      mux_sel = 3'h2;
      done = 1'h1;
    end
  end
  if (~done) begin
    if ((~max_value[3]) & (dimensionality > 4'h3)) begin
      mux_sel = 3'h3;
      done = 1'h1;
    end
  end
  if (~done) begin
    if ((~max_value[4]) & (dimensionality > 4'h4)) begin
      mux_sel = 3'h4;
      done = 1'h1;
    end
  end
  if (~done) begin
    if ((~max_value[5]) & (dimensionality > 4'h5)) begin
      mux_sel = 3'h5;
      done = 1'h1;
    end
  end
end
always_comb begin
  clear[0] = 1'h0;
  if (((mux_sel > 3'h0) | (~done)) & step) begin
    clear[0] = 1'h1;
  end
end
always_comb begin
  inc[0] = 1'h0;
  if ((5'h0 == 5'h0) & step & (dimensionality > 4'h0)) begin
    inc[0] = 1'h1;
  end
  else if ((mux_sel == 3'h0) & step & (dimensionality > 4'h0)) begin
    inc[0] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[0] <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[0] <= 16'h0;
    end
    else if (clear[0]) begin
      dim_counter[0] <= 16'h0;
    end
    else if (inc[0]) begin
      dim_counter[0] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[0] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[0] <= 1'h0;
    end
    else if (clear[0]) begin
      max_value[0] <= 1'h0;
    end
    else if (inc[0]) begin
      max_value[0] <= maxed_value;
    end
  end
end
always_comb begin
  clear[1] = 1'h0;
  if (((mux_sel > 3'h1) | (~done)) & step) begin
    clear[1] = 1'h1;
  end
end
always_comb begin
  inc[1] = 1'h0;
  if ((5'h1 == 5'h0) & step & (dimensionality > 4'h1)) begin
    inc[1] = 1'h1;
  end
  else if ((mux_sel == 3'h1) & step & (dimensionality > 4'h1)) begin
    inc[1] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[1] <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[1] <= 16'h0;
    end
    else if (clear[1]) begin
      dim_counter[1] <= 16'h0;
    end
    else if (inc[1]) begin
      dim_counter[1] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[1] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[1] <= 1'h0;
    end
    else if (clear[1]) begin
      max_value[1] <= 1'h0;
    end
    else if (inc[1]) begin
      max_value[1] <= maxed_value;
    end
  end
end
always_comb begin
  clear[2] = 1'h0;
  if (((mux_sel > 3'h2) | (~done)) & step) begin
    clear[2] = 1'h1;
  end
end
always_comb begin
  inc[2] = 1'h0;
  if ((5'h2 == 5'h0) & step & (dimensionality > 4'h2)) begin
    inc[2] = 1'h1;
  end
  else if ((mux_sel == 3'h2) & step & (dimensionality > 4'h2)) begin
    inc[2] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[2] <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[2] <= 16'h0;
    end
    else if (clear[2]) begin
      dim_counter[2] <= 16'h0;
    end
    else if (inc[2]) begin
      dim_counter[2] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[2] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[2] <= 1'h0;
    end
    else if (clear[2]) begin
      max_value[2] <= 1'h0;
    end
    else if (inc[2]) begin
      max_value[2] <= maxed_value;
    end
  end
end
always_comb begin
  clear[3] = 1'h0;
  if (((mux_sel > 3'h3) | (~done)) & step) begin
    clear[3] = 1'h1;
  end
end
always_comb begin
  inc[3] = 1'h0;
  if ((5'h3 == 5'h0) & step & (dimensionality > 4'h3)) begin
    inc[3] = 1'h1;
  end
  else if ((mux_sel == 3'h3) & step & (dimensionality > 4'h3)) begin
    inc[3] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[3] <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[3] <= 16'h0;
    end
    else if (clear[3]) begin
      dim_counter[3] <= 16'h0;
    end
    else if (inc[3]) begin
      dim_counter[3] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[3] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[3] <= 1'h0;
    end
    else if (clear[3]) begin
      max_value[3] <= 1'h0;
    end
    else if (inc[3]) begin
      max_value[3] <= maxed_value;
    end
  end
end
always_comb begin
  clear[4] = 1'h0;
  if (((mux_sel > 3'h4) | (~done)) & step) begin
    clear[4] = 1'h1;
  end
end
always_comb begin
  inc[4] = 1'h0;
  if ((5'h4 == 5'h0) & step & (dimensionality > 4'h4)) begin
    inc[4] = 1'h1;
  end
  else if ((mux_sel == 3'h4) & step & (dimensionality > 4'h4)) begin
    inc[4] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[4] <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[4] <= 16'h0;
    end
    else if (clear[4]) begin
      dim_counter[4] <= 16'h0;
    end
    else if (inc[4]) begin
      dim_counter[4] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[4] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[4] <= 1'h0;
    end
    else if (clear[4]) begin
      max_value[4] <= 1'h0;
    end
    else if (inc[4]) begin
      max_value[4] <= maxed_value;
    end
  end
end
always_comb begin
  clear[5] = 1'h0;
  if (((mux_sel > 3'h5) | (~done)) & step) begin
    clear[5] = 1'h1;
  end
end
always_comb begin
  inc[5] = 1'h0;
  if ((5'h5 == 5'h0) & step & (dimensionality > 4'h5)) begin
    inc[5] = 1'h1;
  end
  else if ((mux_sel == 3'h5) & step & (dimensionality > 4'h5)) begin
    inc[5] = 1'h1;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    dim_counter[5] <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      dim_counter[5] <= 16'h0;
    end
    else if (clear[5]) begin
      dim_counter[5] <= 16'h0;
    end
    else if (inc[5]) begin
      dim_counter[5] <= inced_cnt;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    max_value[5] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      max_value[5] <= 1'h0;
    end
    else if (clear[5]) begin
      max_value[5] <= 1'h0;
    end
    else if (inc[5]) begin
      max_value[5] <= maxed_value;
    end
  end
end
assign restart = step & (~done);
endmodule   // for_loop_6_16

module reg_fifo_d_4_w_1 #(
  parameter data_width = 16'h10
)
(
  input logic clk,
  input logic clk_en,
  input logic [0:0] [data_width-1:0] data_in,
  input logic flush,
  input logic [2:0] num_load,
  input logic [3:0][0:0] [data_width-1:0] parallel_in,
  input logic parallel_load,
  input logic parallel_read,
  input logic pop,
  input logic push,
  input logic rst_n,
  output logic [0:0] [data_width-1:0] data_out,
  output logic empty,
  output logic full,
  output logic [3:0][0:0] [data_width-1:0] parallel_out,
  output logic [1:0] rd_ptr_out,
  output logic valid
);

logic [2:0] num_items;
logic passthru;
logic [1:0] rd_ptr;
logic read;
logic [3:0][0:0][data_width-1:0] reg_array;
logic [1:0] wr_ptr;
logic write;
assign rd_ptr_out = rd_ptr;
assign full = num_items == 3'h4;
assign empty = num_items == 3'h0;
assign read = pop & (~passthru) & (~empty);
assign passthru = pop & push & empty;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    num_items <= 3'h0;
  end
  else if (flush) begin
    num_items <= 3'h0;
  end
  else if (clk_en) begin
    if (parallel_load) begin
      if (num_load == 3'h0) begin
        num_items <= 3'(push);
      end
      else num_items <= num_load;
    end
    else if (parallel_read) begin
      if (push) begin
        num_items <= 3'h1;
      end
      else num_items <= 3'h0;
    end
    else if (write & (~read)) begin
      num_items <= num_items + 3'h1;
    end
    else if ((~write) & read) begin
      num_items <= num_items - 3'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    reg_array <= 64'h0;
  end
  else if (flush) begin
    reg_array <= 64'h0;
  end
  else if (clk_en) begin
    if (parallel_load) begin
      reg_array <= parallel_in;
    end
    else if (write) begin
      if (parallel_read) begin
        reg_array[0] <= data_in;
      end
      else reg_array[wr_ptr] <= data_in;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    wr_ptr <= 2'h0;
  end
  else if (flush) begin
    wr_ptr <= 2'h0;
  end
  else if (clk_en) begin
    if (parallel_load) begin
      wr_ptr <= num_load[1:0];
    end
    else if (parallel_read) begin
      if (push) begin
        wr_ptr <= 2'h1;
      end
      else wr_ptr <= 2'h0;
    end
    else if (write) begin
      wr_ptr <= wr_ptr + 2'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    rd_ptr <= 2'h0;
  end
  else if (flush) begin
    rd_ptr <= 2'h0;
  end
  else if (clk_en) begin
    if (parallel_load | parallel_read) begin
      rd_ptr <= 2'h0;
    end
    else if (read) begin
      rd_ptr <= rd_ptr + 2'h1;
    end
  end
end
assign parallel_out = reg_array;
assign write = push & (~passthru) & ((~full) | pop | parallel_read);
always_comb begin
  if (passthru) begin
    data_out = data_in;
  end
  else data_out = reg_array[rd_ptr];
end
always_comb begin
  valid = pop & ((~empty) | passthru);
end
endmodule   // reg_fifo_d_4_w_1

module reg_fifo_d_4_w_1_unq0 #(
  parameter data_width = 16'h10
)
(
  input logic clk,
  input logic clk_en,
  input logic [0:0] [data_width-1:0] data_in,
  input logic flush,
  input logic [2:0] num_load,
  input logic [3:0][0:0] [data_width-1:0] parallel_in,
  input logic parallel_load,
  input logic parallel_read,
  input logic pop,
  input logic push,
  input logic rst_n,
  output logic [0:0] [data_width-1:0] data_out,
  output logic empty,
  output logic full,
  output logic [3:0][0:0] [data_width-1:0] parallel_out,
  output logic valid
);

logic [2:0] num_items;
logic passthru;
logic [1:0] rd_ptr;
logic read;
logic [3:0][0:0][data_width-1:0] reg_array;
logic [1:0] wr_ptr;
logic write;
assign full = num_items == 3'h4;
assign empty = num_items == 3'h0;
assign read = pop & (~passthru) & (~empty);
assign passthru = pop & push & empty;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    num_items <= 3'h0;
  end
  else if (flush) begin
    num_items <= 3'h0;
  end
  else if (clk_en) begin
    if (parallel_load) begin
      if (num_load == 3'h0) begin
        num_items <= 3'(push);
      end
      else num_items <= num_load;
    end
    else if (parallel_read) begin
      if (push) begin
        num_items <= 3'h1;
      end
      else num_items <= 3'h0;
    end
    else if (write & (~read)) begin
      num_items <= num_items + 3'h1;
    end
    else if ((~write) & read) begin
      num_items <= num_items - 3'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    reg_array <= 64'h0;
  end
  else if (flush) begin
    reg_array <= 64'h0;
  end
  else if (clk_en) begin
    if (parallel_load) begin
      reg_array <= parallel_in;
    end
    else if (write) begin
      if (parallel_read) begin
        reg_array[0] <= data_in;
      end
      else reg_array[wr_ptr] <= data_in;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    wr_ptr <= 2'h0;
  end
  else if (flush) begin
    wr_ptr <= 2'h0;
  end
  else if (clk_en) begin
    if (parallel_load) begin
      wr_ptr <= num_load[1:0];
    end
    else if (parallel_read) begin
      if (push) begin
        wr_ptr <= 2'h1;
      end
      else wr_ptr <= 2'h0;
    end
    else if (write) begin
      wr_ptr <= wr_ptr + 2'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    rd_ptr <= 2'h0;
  end
  else if (flush) begin
    rd_ptr <= 2'h0;
  end
  else if (clk_en) begin
    if (parallel_load | parallel_read) begin
      rd_ptr <= 2'h0;
    end
    else if (read) begin
      rd_ptr <= rd_ptr + 2'h1;
    end
  end
end
assign parallel_out = reg_array;
assign write = push & (~passthru) & ((~full) | pop | parallel_read);
always_comb begin
  if (passthru) begin
    data_out = data_in;
  end
  else data_out = reg_array[rd_ptr];
end
always_comb begin
  valid = pop & ((~empty) | passthru);
end
endmodule   // reg_fifo_d_4_w_1_unq0

module sched_gen_6_16 (
  input logic clk,
  input logic clk_en,
  input logic [15:0] cycle_count,
  input logic enable,
  input logic finished,
  input logic flush,
  input logic [2:0] mux_sel,
  input logic rst_n,
  input logic [15:0] sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] sched_addr_gen_strides,
  output logic valid_output
);

logic [15:0] addr_out;
logic valid_gate;
logic valid_gate_inv;
logic valid_out;
assign valid_gate = ~valid_gate_inv;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    valid_gate_inv <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      valid_gate_inv <= 1'h0;
    end
    else if (finished) begin
      valid_gate_inv <= 1'h1;
    end
  end
end
always_comb begin
  valid_out = (cycle_count == addr_out) & valid_gate & enable;
end
always_comb begin
  valid_output = valid_out;
end
addr_gen_6_16 sched_addr_gen (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(mux_sel),
  .restart(1'h0),
  .rst_n(rst_n),
  .starting_addr(sched_addr_gen_starting_addr),
  .step(valid_out),
  .strides(sched_addr_gen_strides),
  .addr_out(addr_out)
);

endmodule   // sched_gen_6_16

module sram_stub (
  input logic [8:0] addr,
  input logic cen,
  input logic clk,
  input logic clk_en,
  input logic [3:0] [15:0] data_in,
  input logic flush,
  input logic wen,
  output logic [3:0] [15:0] data_out
);

logic [511:0][3:0][15:0] data_array;

always_ff @(posedge clk) begin
  if (clk_en) begin
    if (cen & wen) begin
      data_array[addr] <= data_in;
    end
  end
end

always_ff @(posedge clk) begin
  if (clk_en) begin
    if (cen & (~wen)) begin
      data_out <= data_array[addr];
    end
  end
end
endmodule   // sram_stub

module storage_config_seq (
  input logic clk,
  input logic clk_en,
  input logic [7:0] config_addr_in,
  input logic [15:0] config_data_in,
  input logic [1:0] config_en,
  input logic config_rd,
  input logic config_wr,
  input logic flush,
  input logic [0:0][3:0] [15:0] rd_data_stg,
  input logic rst_n,
  output logic [8:0] addr_out,
  output logic [1:0] [15:0] rd_data_out,
  output logic ren_out,
  output logic wen_out,
  output logic [3:0] [15:0] wr_data
);

logic [1:0] cnt;
logic [2:0][15:0] data_wr_reg;
logic [1:0] rd_cnt;
logic [1:0] reduce_en;
logic set_to_addr;
assign reduce_en[0] = |config_en[0];
assign reduce_en[1] = |config_en[1];
always_comb begin
  set_to_addr = 1'h0;
  for (int unsigned i = 0; i < 2; i += 1) begin
      if (reduce_en[1'(i)]) begin
        set_to_addr = 1'(i);
      end
    end
end
assign addr_out = {set_to_addr, config_addr_in};

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    cnt <= 2'h0;
  end
  else if (flush) begin
    cnt <= 2'h0;
  end
  else if (clk_en) begin
    if ((config_wr | config_rd) & (|config_en)) begin
      cnt <= cnt + 2'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    rd_cnt <= 2'h0;
  end
  else if (flush) begin
    rd_cnt <= 2'h0;
  end
  else if (clk_en) begin
    rd_cnt <= cnt;
  end
end
assign rd_data_out[0] = rd_data_stg[0][rd_cnt];
assign rd_data_out[1] = rd_data_stg[0][rd_cnt];

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    data_wr_reg <= 48'h0;
  end
  else if (flush) begin
    data_wr_reg <= 48'h0;
  end
  else if (clk_en) begin
    if (config_wr & (cnt < 2'h3)) begin
      data_wr_reg[cnt] <= config_data_in;
    end
  end
end
assign wr_data[0] = data_wr_reg[0];
assign wr_data[1] = data_wr_reg[1];
assign wr_data[2] = data_wr_reg[2];
assign wr_data[3] = config_data_in;
assign wen_out = config_wr & (cnt == 2'h3);
assign ren_out = config_rd;
endmodule   // storage_config_seq

module strg_fifo (
  input logic clk,
  input logic clk_en,
  input logic [0:0][3:0] [15:0] data_from_strg,
  input logic [15:0] data_in,
  input logic [15:0] fifo_depth,
  input logic flush,
  input logic pop,
  input logic push,
  input logic rst_n,
  output logic [0:0] [8:0] addr_out,
  output logic [15:0] data_out,
  output logic [0:0][3:0] [15:0] data_to_strg,
  output logic empty,
  output logic full,
  output logic ren_to_strg,
  output logic valid_out,
  output logic wen_to_strg
);

logic [15:0] back_data_in;
logic [15:0] back_data_out;
logic back_empty;
logic back_full;
logic [2:0] back_num_load;
logic [2:0] back_occ;
logic [3:0][0:0][15:0] back_par_in;
logic back_pl;
logic back_pop;
logic back_push;
logic [0:0][15:0] back_rf_data_in;
logic [0:0][15:0] back_rf_data_out;
logic back_rf_parallel_load;
logic back_valid;
logic curr_bank_rd;
logic curr_bank_wr;
logic [3:0][15:0] front_combined;
logic [15:0] front_data_out;
logic front_empty;
logic front_full;
logic [2:0] front_occ;
logic [3:0][0:0][15:0] front_par_out;
logic front_par_read;
logic front_pop;
logic front_push;
logic [1:0] front_rd_ptr;
logic [0:0][15:0] front_rf_data_in;
logic [0:0][15:0] front_rf_data_out;
logic front_valid;
logic fw_is_1;
logic [15:0] num_items;
logic [15:0] num_words_mem;
logic prev_bank_rd;
logic queued_write;
logic [0:0][8:0] ren_addr;
logic ren_delay;
logic [0:0][8:0] wen_addr;
logic [0:0][3:0][15:0] write_queue;
assign curr_bank_wr = 1'h0;
assign curr_bank_rd = 1'h0;
assign front_push = push & ((~full) | pop);
assign front_rf_data_in[0] = data_in;
assign front_data_out = front_rf_data_out[0];
assign fw_is_1 = 1'h0;
assign back_pop = pop & ((~empty) | push);
assign back_rf_parallel_load = back_pl & (|back_num_load);
assign back_rf_data_in[0] = back_data_in;
assign back_data_out = back_rf_data_out[0];
always_comb begin
  wen_to_strg = ((~ren_to_strg) | 1'h0) & (queued_write | ((front_occ == 3'h4) & push &
      (~front_pop) & (curr_bank_wr == 1'h0)));
end
always_comb begin
  ren_to_strg = ((back_occ == 3'h1) | fw_is_1) & (curr_bank_rd == 1'h0) & (pop | ((back_occ ==
      3'h0) & (back_num_load == 3'h0))) & ((num_words_mem > 16'h1) | ((num_words_mem
      == 16'h1) & (~back_pl)));
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    ren_delay <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      ren_delay <= 1'h0;
    end
    else ren_delay <= |ren_to_strg;
  end
end
assign back_pl = ren_delay;
assign front_combined[0] = front_par_out[front_rd_ptr + 2'h0];
assign front_combined[1] = front_par_out[front_rd_ptr + 2'h1];
assign front_combined[2] = front_par_out[front_rd_ptr + 2'h2];
assign front_combined[3] = front_par_out[front_rd_ptr + 2'h3];
assign data_to_strg[0] = queued_write ? write_queue[0]: front_combined;
assign back_data_in = front_data_out;
assign back_push = front_valid;
always_comb begin
  front_pop = ((num_words_mem == 16'h0) | ((num_words_mem == 16'h1) & back_pl)) & ((~back_pl)
      | (back_pl & (back_num_load == 3'h0))) & ((~(back_occ == 3'h4)) | pop) &
      ((~(front_occ == 3'h0)) | push);
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    write_queue[0] <= 64'h0;
    queued_write <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      write_queue[0] <= 64'h0;
      queued_write <= 1'h0;
    end
    else if (front_par_read & (~wen_to_strg) & (curr_bank_wr == 1'h0)) begin
      write_queue[0] <= front_combined;
      queued_write <= 1'h1;
    end
    else if (wen_to_strg) begin
      queued_write <= 1'h0;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    num_words_mem <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      num_words_mem <= 16'h0;
    end
    else if ((~back_pl) & front_par_read) begin
      num_words_mem <= num_words_mem + 16'h1;
    end
    else if (back_pl & (~front_par_read)) begin
      num_words_mem <= num_words_mem - 16'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    front_occ <= 3'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      front_occ <= 3'h0;
    end
    else if (front_par_read) begin
      if (front_push) begin
        front_occ <= 3'h1;
      end
      else front_occ <= 3'h0;
    end
    else if (front_push & (~front_pop)) begin
      front_occ <= front_occ + 3'h1;
    end
    else if ((~front_push) & front_pop) begin
      front_occ <= front_occ - 3'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    back_occ <= 3'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      back_occ <= 3'h0;
    end
    else if (back_pl) begin
      if (back_num_load == 3'h0) begin
        back_occ <= 3'(back_push);
      end
      else back_occ <= back_num_load;
    end
    else if (back_push & (~back_pop)) begin
      back_occ <= back_occ + 3'h1;
    end
    else if ((~back_push) & back_pop) begin
      back_occ <= back_occ - 3'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    prev_bank_rd <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      prev_bank_rd <= 1'h0;
    end
    else prev_bank_rd <= curr_bank_rd;
  end
end
assign back_par_in[0] = (back_num_load == 3'h4) ? data_from_strg[prev_bank_rd][0]:
    data_from_strg[prev_bank_rd][1];
assign back_par_in[1] = (back_num_load == 3'h4) ? data_from_strg[prev_bank_rd][1]:
    data_from_strg[prev_bank_rd][2];
assign back_par_in[2] = (back_num_load == 3'h4) ? data_from_strg[prev_bank_rd][2]:
    data_from_strg[prev_bank_rd][3];
assign back_par_in[3] = (back_num_load == 3'h4) ? data_from_strg[prev_bank_rd][3]: 16'h0;
always_comb begin
  front_par_read = (front_occ == 3'h4) & push & (~front_pop);
end
always_comb begin
  if (back_pl) begin
    back_num_load = pop ? 3'h3: 3'h4;
  end
  else back_num_load = 3'h0;
end
assign data_out = back_pl ? data_from_strg[prev_bank_rd][0]: back_data_out;
assign valid_out = back_pl ? pop: back_valid;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    wen_addr[0] <= 9'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      wen_addr[0] <= 9'h0;
    end
    else if (wen_to_strg) begin
      wen_addr[0] <= wen_addr[0] + 9'h1;
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    ren_addr[0] <= 9'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      ren_addr[0] <= 9'h0;
    end
    else if (ren_to_strg) begin
      ren_addr[0] <= ren_addr[0] + 9'h1;
    end
  end
end
assign addr_out[0] = wen_to_strg ? wen_addr[0]: ren_addr[0];
always_comb begin
  num_items = 16'(num_words_mem * 16'h4) + 16'(front_occ) + 16'(back_occ);
end
assign empty = num_items == 16'h0;
assign full = fifo_depth == num_items;
reg_fifo_d_4_w_1 #(
  .data_width(16'h10))
front_rf (
  .clk(clk),
  .clk_en(clk_en),
  .data_in(front_rf_data_in),
  .flush(flush),
  .num_load(3'h0),
  .parallel_in(64'h0),
  .parallel_load(1'h0),
  .parallel_read(front_par_read),
  .pop(front_pop),
  .push(front_push),
  .rst_n(rst_n),
  .data_out(front_rf_data_out),
  .empty(front_empty),
  .full(front_full),
  .parallel_out(front_par_out),
  .rd_ptr_out(front_rd_ptr),
  .valid(front_valid)
);

reg_fifo_d_4_w_1_unq0 #(
  .data_width(16'h10))
back_rf (
  .clk(clk),
  .clk_en(clk_en),
  .data_in(back_rf_data_in),
  .flush(flush),
  .num_load(back_num_load),
  .parallel_in(back_par_in),
  .parallel_load(back_rf_parallel_load),
  .parallel_read(1'h0),
  .pop(back_pop),
  .push(back_push),
  .rst_n(rst_n),
  .data_out(back_rf_data_out),
  .empty(back_empty),
  .full(back_full),
  .valid(back_valid)
);

endmodule   // strg_fifo

module strg_ram (
  input logic clk,
  input logic clk_en,
  input logic [0:0][3:0] [15:0] data_from_strg,
  input logic [15:0] data_in,
  input logic flush,
  input logic [15:0] rd_addr_in,
  input logic ren,
  input logic rst_n,
  input logic wen,
  input logic [15:0] wr_addr_in,
  output logic [0:0] [8:0] addr_out,
  output logic [15:0] data_out,
  output logic [0:0][3:0] [15:0] data_to_strg,
  output logic ready,
  output logic ren_to_strg,
  output logic valid_out,
  output logic wen_to_strg
);

typedef enum logic[1:0] {
  IDLE = 2'h0,
  MODIFY = 2'h1,
  READ = 2'h2,
  _DEFAULT = 2'h3
} r_w_seq_state;
logic [15:0] addr_to_write;
logic [3:0][15:0] data_combined;
logic [15:0] data_to_write;
r_w_seq_state r_w_seq_current_state;
r_w_seq_state r_w_seq_next_state;
logic [15:0] rd_addr;
logic rd_bank;
logic rd_valid;
logic read_gate;
logic [15:0] wr_addr;
logic write_gate;
assign wr_addr = wr_addr_in;
assign rd_addr = wr_addr_in;
assign rd_bank = 1'h0;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    rd_valid <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      rd_valid <= 1'h0;
    end
    else rd_valid <= ren & (~wen);
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    data_to_write <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      data_to_write <= 16'h0;
    end
    else data_to_write <= data_in;
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    addr_to_write <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      addr_to_write <= 16'h0;
    end
    else addr_to_write <= wr_addr;
  end
end
assign data_to_strg[0] = data_combined;
assign ren_to_strg = (wen | ren) & read_gate;
assign wen_to_strg = write_gate;
always_comb begin
  addr_out[0] = rd_addr[10:2];
  if (wen & (~write_gate)) begin
    addr_out[0] = wr_addr[10:2];
  end
  else if (write_gate) begin
    addr_out[0] = addr_to_write[10:2];
  end
end
always_comb begin
  if (addr_to_write[1:0] == 2'h0) begin
    data_combined[0] = data_to_write;
  end
  else data_combined[0] = data_from_strg[rd_bank][0];
end
always_comb begin
  if (addr_to_write[1:0] == 2'h1) begin
    data_combined[1] = data_to_write;
  end
  else data_combined[1] = data_from_strg[rd_bank][1];
end
always_comb begin
  if (addr_to_write[1:0] == 2'h2) begin
    data_combined[2] = data_to_write;
  end
  else data_combined[2] = data_from_strg[rd_bank][2];
end
always_comb begin
  if (addr_to_write[1:0] == 2'h3) begin
    data_combined[3] = data_to_write;
  end
  else data_combined[3] = data_from_strg[rd_bank][3];
end

always_ff @(posedge clk, negedge rst_n) begin
  if (!rst_n) begin
    r_w_seq_current_state <= IDLE;
  end
  else r_w_seq_current_state <= r_w_seq_next_state;
end
always_comb begin
  r_w_seq_next_state = r_w_seq_current_state;
  unique case (r_w_seq_current_state)
    IDLE: begin
        if ((~wen) & (~ren)) begin
          r_w_seq_next_state = IDLE;
        end
        else if (wen) begin
          r_w_seq_next_state = MODIFY;
        end
        else if (ren & (~wen)) begin
          r_w_seq_next_state = READ;
        end
      end
    MODIFY: begin
        if (1'h1) begin
          r_w_seq_next_state = IDLE;
        end
      end
    READ: begin
        if ((~wen) & (~ren)) begin
          r_w_seq_next_state = IDLE;
        end
        else if (wen) begin
          r_w_seq_next_state = MODIFY;
        end
        else if (ren & (~wen)) begin
          r_w_seq_next_state = READ;
        end
      end
    _DEFAULT: begin
        if (1'h1) begin
          r_w_seq_next_state = _DEFAULT;
        end
      end
  endcase
end
always_comb begin
  unique case (r_w_seq_current_state)
    IDLE: begin :r_w_seq_IDLE_Output
        data_out = 16'h0;
        read_gate = 1'h1;
        ready = 1'h1;
        valid_out = 1'h0;
        write_gate = 1'h0;
      end :r_w_seq_IDLE_Output
    MODIFY: begin :r_w_seq_MODIFY_Output
        data_out = 16'h0;
        read_gate = 1'h0;
        ready = 1'h0;
        valid_out = 1'h0;
        write_gate = 1'h1;
      end :r_w_seq_MODIFY_Output
    READ: begin :r_w_seq_READ_Output
        data_out = data_from_strg[rd_bank][addr_to_write[1:0]];
        read_gate = 1'h1;
        ready = 1'h1;
        valid_out = 1'h1;
        write_gate = 1'h0;
      end :r_w_seq_READ_Output
    _DEFAULT: begin :r_w_seq__DEFAULT_Output
        data_out = 16'h0;
        read_gate = 1'h0;
        ready = 1'h0;
        valid_out = 1'h0;
        write_gate = 1'h0;
      end :r_w_seq__DEFAULT_Output
  endcase
end
endmodule   // strg_ram

module strg_ub_agg_only (
  input logic [1:0] agg_read,
  input logic [3:0] agg_read_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] agg_read_addr_gen_0_strides,
  input logic [3:0] agg_read_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] agg_read_addr_gen_1_strides,
  input logic [3:0] agg_write_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] agg_write_addr_gen_0_strides,
  input logic [3:0] agg_write_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] agg_write_addr_gen_1_strides,
  input logic agg_write_sched_gen_0_enable,
  input logic [15:0] agg_write_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] agg_write_sched_gen_0_sched_addr_gen_strides,
  input logic agg_write_sched_gen_1_enable,
  input logic [15:0] agg_write_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] agg_write_sched_gen_1_sched_addr_gen_strides,
  input logic clk,
  input logic clk_en,
  input logic [15:0] cycle_count,
  input logic [1:0] [15:0] data_in,
  input logic [1:0] [2:0] floop_mux_sel,
  input logic [1:0] floop_restart,
  input logic flush,
  input logic [3:0] loops_in2buf_0_dimensionality,
  input logic [5:0] [15:0] loops_in2buf_0_ranges,
  input logic [3:0] loops_in2buf_1_dimensionality,
  input logic [5:0] [15:0] loops_in2buf_1_ranges,
  input logic rst_n,
  output logic [1:0][3:0] [15:0] agg_data_out
);

logic [1:0][3:0][3:0][15:0] agg;
logic [1:0][1:0] agg_read_addr;
logic [3:0] agg_read_addr_gen_0_addr_out;
logic [2:0] agg_read_addr_gen_0_mux_sel;
logic agg_read_addr_gen_0_restart;
logic agg_read_addr_gen_0_step;
logic [3:0] agg_read_addr_gen_1_addr_out;
logic [2:0] agg_read_addr_gen_1_mux_sel;
logic agg_read_addr_gen_1_restart;
logic agg_read_addr_gen_1_step;
logic [1:0][7:0] agg_read_addr_gen_out;
logic [1:0] agg_write;
logic [1:0][3:0] agg_write_addr;
logic [3:0] agg_write_addr_gen_0_addr_out;
logic agg_write_addr_gen_0_step;
logic [3:0] agg_write_addr_gen_1_addr_out;
logic agg_write_addr_gen_1_step;
logic agg_write_sched_gen_0_valid_output;
logic agg_write_sched_gen_1_valid_output;
logic [2:0] loops_in2buf_0_mux_sel_out;
logic loops_in2buf_0_restart;
logic loops_in2buf_0_step;
logic [2:0] loops_in2buf_1_mux_sel_out;
logic loops_in2buf_1_restart;
logic loops_in2buf_1_step;
assign loops_in2buf_0_step = agg_write[0];
assign agg_write_addr_gen_0_step = agg_write[0];
assign agg_write_addr[0] = agg_write_addr_gen_0_addr_out;
assign agg_write[0] = agg_write_sched_gen_0_valid_output;

always_ff @(posedge clk) begin
  if (clk_en) begin
    if (agg_write[0]) begin
      agg[0][agg_write_addr[0][3:2]][agg_write_addr[0][1:0]] <= data_in[0];
    end
  end
end
assign agg_read_addr_gen_0_step = agg_read[0];
assign agg_read_addr_gen_0_restart = floop_restart[0];
assign agg_read_addr_gen_0_mux_sel = floop_mux_sel[0];
assign agg_read_addr_gen_out[0][3:0] = agg_read_addr_gen_0_addr_out;
assign agg_read_addr_gen_out[0][7:4] = 4'h0;
assign agg_read_addr[0] = agg_read_addr_gen_out[0][1:0];
always_comb begin
  agg_data_out[0] = agg[0][agg_read_addr[0]];
end
assign loops_in2buf_1_step = agg_write[1];
assign agg_write_addr_gen_1_step = agg_write[1];
assign agg_write_addr[1] = agg_write_addr_gen_1_addr_out;
assign agg_write[1] = agg_write_sched_gen_1_valid_output;

always_ff @(posedge clk) begin
  if (clk_en) begin
    if (agg_write[1]) begin
      agg[1][agg_write_addr[1][3:2]][agg_write_addr[1][1:0]] <= data_in[1];
    end
  end
end
assign agg_read_addr_gen_1_step = agg_read[1];
assign agg_read_addr_gen_1_restart = floop_restart[1];
assign agg_read_addr_gen_1_mux_sel = floop_mux_sel[1];
assign agg_read_addr_gen_out[1][3:0] = agg_read_addr_gen_1_addr_out;
assign agg_read_addr_gen_out[1][7:4] = 4'h0;
assign agg_read_addr[1] = agg_read_addr_gen_out[1][1:0];
always_comb begin
  agg_data_out[1] = agg[1][agg_read_addr[1]];
end
for_loop_6_16 #(
  .CONFIG_WIDTH(5'h10),
  .ITERATOR_SUPPORT(4'h6))
loops_in2buf_0 (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_in2buf_0_dimensionality),
  .flush(flush),
  .ranges(loops_in2buf_0_ranges),
  .rst_n(rst_n),
  .step(loops_in2buf_0_step),
  .mux_sel_out(loops_in2buf_0_mux_sel_out),
  .restart(loops_in2buf_0_restart)
);

addr_gen_6_4 agg_write_addr_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(loops_in2buf_0_mux_sel_out),
  .restart(loops_in2buf_0_restart),
  .rst_n(rst_n),
  .starting_addr(agg_write_addr_gen_0_starting_addr),
  .step(agg_write_addr_gen_0_step),
  .strides(agg_write_addr_gen_0_strides),
  .addr_out(agg_write_addr_gen_0_addr_out)
);

sched_gen_6_16 agg_write_sched_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(agg_write_sched_gen_0_enable),
  .finished(loops_in2buf_0_restart),
  .flush(flush),
  .mux_sel(loops_in2buf_0_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(agg_write_sched_gen_0_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides(agg_write_sched_gen_0_sched_addr_gen_strides),
  .valid_output(agg_write_sched_gen_0_valid_output)
);

addr_gen_6_4 agg_read_addr_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(agg_read_addr_gen_0_mux_sel),
  .restart(agg_read_addr_gen_0_restart),
  .rst_n(rst_n),
  .starting_addr(agg_read_addr_gen_0_starting_addr),
  .step(agg_read_addr_gen_0_step),
  .strides(agg_read_addr_gen_0_strides),
  .addr_out(agg_read_addr_gen_0_addr_out)
);

for_loop_6_16 #(
  .CONFIG_WIDTH(5'h10),
  .ITERATOR_SUPPORT(4'h6))
loops_in2buf_1 (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_in2buf_1_dimensionality),
  .flush(flush),
  .ranges(loops_in2buf_1_ranges),
  .rst_n(rst_n),
  .step(loops_in2buf_1_step),
  .mux_sel_out(loops_in2buf_1_mux_sel_out),
  .restart(loops_in2buf_1_restart)
);

addr_gen_6_4 agg_write_addr_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(loops_in2buf_1_mux_sel_out),
  .restart(loops_in2buf_1_restart),
  .rst_n(rst_n),
  .starting_addr(agg_write_addr_gen_1_starting_addr),
  .step(agg_write_addr_gen_1_step),
  .strides(agg_write_addr_gen_1_strides),
  .addr_out(agg_write_addr_gen_1_addr_out)
);

sched_gen_6_16 agg_write_sched_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(agg_write_sched_gen_1_enable),
  .finished(loops_in2buf_1_restart),
  .flush(flush),
  .mux_sel(loops_in2buf_1_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(agg_write_sched_gen_1_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides(agg_write_sched_gen_1_sched_addr_gen_strides),
  .valid_output(agg_write_sched_gen_1_valid_output)
);

addr_gen_6_4 agg_read_addr_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(agg_read_addr_gen_1_mux_sel),
  .restart(agg_read_addr_gen_1_restart),
  .rst_n(rst_n),
  .starting_addr(agg_read_addr_gen_1_starting_addr),
  .step(agg_read_addr_gen_1_step),
  .strides(agg_read_addr_gen_1_strides),
  .addr_out(agg_read_addr_gen_1_addr_out)
);

endmodule   // strg_ub_agg_only

module strg_ub_agg_sram_shared (
  input logic agg_read_sched_gen_0_enable,
  input logic [15:0] agg_read_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] agg_read_sched_gen_0_sched_addr_gen_strides,
  input logic agg_read_sched_gen_1_enable,
  input logic [15:0] agg_read_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] agg_read_sched_gen_1_sched_addr_gen_strides,
  input logic clk,
  input logic clk_en,
  input logic [15:0] cycle_count,
  input logic flush,
  input logic [3:0] loops_in2buf_autovec_write_0_dimensionality,
  input logic [5:0] [15:0] loops_in2buf_autovec_write_0_ranges,
  input logic [3:0] loops_in2buf_autovec_write_1_dimensionality,
  input logic [5:0] [15:0] loops_in2buf_autovec_write_1_ranges,
  input logic rst_n,
  output logic [1:0] agg_read_out,
  output logic [1:0] [2:0] floop_mux_sel,
  output logic [1:0] floop_restart
);

logic [1:0] agg_read;
logic agg_read_sched_gen_0_valid_output;
logic agg_read_sched_gen_1_valid_output;
logic [2:0] loops_in2buf_autovec_write_0_mux_sel_out;
logic loops_in2buf_autovec_write_0_restart;
logic loops_in2buf_autovec_write_0_step;
logic [2:0] loops_in2buf_autovec_write_1_mux_sel_out;
logic loops_in2buf_autovec_write_1_restart;
logic loops_in2buf_autovec_write_1_step;
assign agg_read_out = agg_read;
assign loops_in2buf_autovec_write_0_step = agg_read[0];
assign floop_mux_sel[0] = loops_in2buf_autovec_write_0_mux_sel_out;
assign floop_restart[0] = loops_in2buf_autovec_write_0_restart;
assign agg_read[0] = agg_read_sched_gen_0_valid_output;
assign loops_in2buf_autovec_write_1_step = agg_read[1];
assign floop_mux_sel[1] = loops_in2buf_autovec_write_1_mux_sel_out;
assign floop_restart[1] = loops_in2buf_autovec_write_1_restart;
assign agg_read[1] = agg_read_sched_gen_1_valid_output;
for_loop_6_16 #(
  .CONFIG_WIDTH(5'h10),
  .ITERATOR_SUPPORT(4'h6))
loops_in2buf_autovec_write_0 (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_in2buf_autovec_write_0_dimensionality),
  .flush(flush),
  .ranges(loops_in2buf_autovec_write_0_ranges),
  .rst_n(rst_n),
  .step(loops_in2buf_autovec_write_0_step),
  .mux_sel_out(loops_in2buf_autovec_write_0_mux_sel_out),
  .restart(loops_in2buf_autovec_write_0_restart)
);

sched_gen_6_16 agg_read_sched_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(agg_read_sched_gen_0_enable),
  .finished(loops_in2buf_autovec_write_0_restart),
  .flush(flush),
  .mux_sel(loops_in2buf_autovec_write_0_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(agg_read_sched_gen_0_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides(agg_read_sched_gen_0_sched_addr_gen_strides),
  .valid_output(agg_read_sched_gen_0_valid_output)
);

for_loop_6_16 #(
  .CONFIG_WIDTH(5'h10),
  .ITERATOR_SUPPORT(4'h6))
loops_in2buf_autovec_write_1 (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_in2buf_autovec_write_1_dimensionality),
  .flush(flush),
  .ranges(loops_in2buf_autovec_write_1_ranges),
  .rst_n(rst_n),
  .step(loops_in2buf_autovec_write_1_step),
  .mux_sel_out(loops_in2buf_autovec_write_1_mux_sel_out),
  .restart(loops_in2buf_autovec_write_1_restart)
);

sched_gen_6_16 agg_read_sched_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(agg_read_sched_gen_1_enable),
  .finished(loops_in2buf_autovec_write_1_restart),
  .flush(flush),
  .mux_sel(loops_in2buf_autovec_write_1_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(agg_read_sched_gen_1_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides(agg_read_sched_gen_1_sched_addr_gen_strides),
  .valid_output(agg_read_sched_gen_1_valid_output)
);

endmodule   // strg_ub_agg_sram_shared

module strg_ub_sram_only (
  input logic [1:0][3:0] [15:0] agg_data_out,
  input logic [1:0] agg_read,
  input logic clk,
  input logic clk_en,
  input logic [15:0] cycle_count,
  input logic [1:0] [2:0] floop_mux_sel,
  input logic [1:0] floop_restart,
  input logic flush,
  input logic [8:0] input_addr_gen_0_starting_addr,
  input logic [5:0] [8:0] input_addr_gen_0_strides,
  input logic [8:0] input_addr_gen_1_starting_addr,
  input logic [5:0] [8:0] input_addr_gen_1_strides,
  input logic [1:0] [2:0] loops_sram2tb_mux_sel,
  input logic [1:0] loops_sram2tb_restart,
  input logic [8:0] output_addr_gen_0_starting_addr,
  input logic [5:0] [8:0] output_addr_gen_0_strides,
  input logic [8:0] output_addr_gen_1_starting_addr,
  input logic [5:0] [8:0] output_addr_gen_1_strides,
  input logic rst_n,
  input logic [1:0] t_read,
  output logic [8:0] addr_to_sram,
  output logic cen_to_sram,
  output logic [3:0] [15:0] data_to_sram,
  output logic wen_to_sram
);

logic [8:0] addr;
logic [3:0][15:0] decode_ret_agg_read_agg_data_out;
logic [15:0] decode_ret_agg_read_s_write_addr;
logic [15:0] decode_ret_t_read_s_read_addr;
logic decode_sel_done_agg_read_agg_data_out;
logic decode_sel_done_agg_read_s_write_addr;
logic decode_sel_done_t_read_s_read_addr;
logic [8:0] input_addr_gen_0_addr_out;
logic [2:0] input_addr_gen_0_mux_sel;
logic input_addr_gen_0_restart;
logic input_addr_gen_0_step;
logic [8:0] input_addr_gen_1_addr_out;
logic [2:0] input_addr_gen_1_mux_sel;
logic input_addr_gen_1_restart;
logic input_addr_gen_1_step;
logic [8:0] output_addr_gen_0_addr_out;
logic [2:0] output_addr_gen_0_mux_sel;
logic output_addr_gen_0_restart;
logic output_addr_gen_0_step;
logic [8:0] output_addr_gen_1_addr_out;
logic [2:0] output_addr_gen_1_mux_sel;
logic output_addr_gen_1_restart;
logic output_addr_gen_1_step;
logic read;
logic [1:0][15:0] s_read_addr;
logic [1:0][15:0] s_write_addr;
logic [3:0][15:0] sram_write_data;
logic write;
assign input_addr_gen_0_step = agg_read[0];
assign input_addr_gen_0_restart = floop_restart[0];
assign input_addr_gen_0_mux_sel = floop_mux_sel[0];
assign s_write_addr[0][8:0] = input_addr_gen_0_addr_out;
assign s_write_addr[0][15:9] = 7'h0;
assign input_addr_gen_1_step = agg_read[1];
assign input_addr_gen_1_restart = floop_restart[1];
assign input_addr_gen_1_mux_sel = floop_mux_sel[1];
assign s_write_addr[1][8:0] = input_addr_gen_1_addr_out;
assign s_write_addr[1][15:9] = 7'h0;
assign output_addr_gen_0_step = t_read[0];
assign output_addr_gen_0_restart = loops_sram2tb_restart[0];
assign output_addr_gen_0_mux_sel = loops_sram2tb_mux_sel[0];
assign s_read_addr[0][8:0] = output_addr_gen_0_addr_out;
assign s_read_addr[0][15:9] = 7'h0;
assign output_addr_gen_1_step = t_read[1];
assign output_addr_gen_1_restart = loops_sram2tb_restart[1];
assign output_addr_gen_1_mux_sel = loops_sram2tb_mux_sel[1];
assign s_read_addr[1][8:0] = output_addr_gen_1_addr_out;
assign s_read_addr[1][15:9] = 7'h0;
assign addr_to_sram = addr;
assign data_to_sram = sram_write_data;
assign wen_to_sram = write;
assign cen_to_sram = write | read;
assign write = |agg_read;
assign read = |t_read;
always_comb begin
  decode_sel_done_agg_read_agg_data_out = 1'h0;
  decode_ret_agg_read_agg_data_out = 64'h0;
  for (int unsigned i = 0; i < 2; i += 1) begin
      if ((~decode_sel_done_agg_read_agg_data_out) & agg_read[1'(i)]) begin
        decode_ret_agg_read_agg_data_out = agg_data_out[1'(i)];
        decode_sel_done_agg_read_agg_data_out = 1'h1;
      end
    end
end
assign sram_write_data = decode_ret_agg_read_agg_data_out;
always_comb begin
  decode_sel_done_agg_read_s_write_addr = 1'h0;
  decode_ret_agg_read_s_write_addr = 16'h0;
  for (int unsigned i = 0; i < 2; i += 1) begin
      if ((~decode_sel_done_agg_read_s_write_addr) & agg_read[1'(i)]) begin
        decode_ret_agg_read_s_write_addr = s_write_addr[1'(i)];
        decode_sel_done_agg_read_s_write_addr = 1'h1;
      end
    end
end
always_comb begin
  decode_sel_done_t_read_s_read_addr = 1'h0;
  decode_ret_t_read_s_read_addr = 16'h0;
  for (int unsigned i = 0; i < 2; i += 1) begin
      if ((~decode_sel_done_t_read_s_read_addr) & t_read[1'(i)]) begin
        decode_ret_t_read_s_read_addr = s_read_addr[1'(i)];
        decode_sel_done_t_read_s_read_addr = 1'h1;
      end
    end
end
always_comb begin
  if (write) begin
    addr = decode_ret_agg_read_s_write_addr[8:0];
  end
  else addr = decode_ret_t_read_s_read_addr[8:0];
end
addr_gen_6_9 input_addr_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(input_addr_gen_0_mux_sel),
  .restart(input_addr_gen_0_restart),
  .rst_n(rst_n),
  .starting_addr(input_addr_gen_0_starting_addr),
  .step(input_addr_gen_0_step),
  .strides(input_addr_gen_0_strides),
  .addr_out(input_addr_gen_0_addr_out)
);

addr_gen_6_9 input_addr_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(input_addr_gen_1_mux_sel),
  .restart(input_addr_gen_1_restart),
  .rst_n(rst_n),
  .starting_addr(input_addr_gen_1_starting_addr),
  .step(input_addr_gen_1_step),
  .strides(input_addr_gen_1_strides),
  .addr_out(input_addr_gen_1_addr_out)
);

addr_gen_6_9 output_addr_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(output_addr_gen_0_mux_sel),
  .restart(output_addr_gen_0_restart),
  .rst_n(rst_n),
  .starting_addr(output_addr_gen_0_starting_addr),
  .step(output_addr_gen_0_step),
  .strides(output_addr_gen_0_strides),
  .addr_out(output_addr_gen_0_addr_out)
);

addr_gen_6_9 output_addr_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(output_addr_gen_1_mux_sel),
  .restart(output_addr_gen_1_restart),
  .rst_n(rst_n),
  .starting_addr(output_addr_gen_1_starting_addr),
  .step(output_addr_gen_1_step),
  .strides(output_addr_gen_1_strides),
  .addr_out(output_addr_gen_1_addr_out)
);

endmodule   // strg_ub_sram_only

module strg_ub_sram_tb_shared (
  input logic clk,
  input logic clk_en,
  input logic [15:0] cycle_count,
  input logic flush,
  input logic [3:0] loops_buf2out_autovec_read_0_dimensionality,
  input logic [5:0] [15:0] loops_buf2out_autovec_read_0_ranges,
  input logic [3:0] loops_buf2out_autovec_read_1_dimensionality,
  input logic [5:0] [15:0] loops_buf2out_autovec_read_1_ranges,
  input logic output_sched_gen_0_enable,
  input logic [15:0] output_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] output_sched_gen_0_sched_addr_gen_strides,
  input logic output_sched_gen_1_enable,
  input logic [15:0] output_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] output_sched_gen_1_sched_addr_gen_strides,
  input logic rst_n,
  output logic [1:0] [2:0] loops_sram2tb_mux_sel,
  output logic [1:0] loops_sram2tb_restart,
  output logic [1:0] t_read_out
);

logic [2:0] loops_buf2out_autovec_read_0_mux_sel_out;
logic loops_buf2out_autovec_read_0_restart;
logic loops_buf2out_autovec_read_0_step;
logic [2:0] loops_buf2out_autovec_read_1_mux_sel_out;
logic loops_buf2out_autovec_read_1_restart;
logic loops_buf2out_autovec_read_1_step;
logic output_sched_gen_0_valid_output;
logic output_sched_gen_1_valid_output;
logic [1:0] t_read;
assign t_read_out = t_read;
assign loops_buf2out_autovec_read_0_step = t_read[0];
assign loops_sram2tb_mux_sel[0] = loops_buf2out_autovec_read_0_mux_sel_out;
assign loops_sram2tb_restart[0] = loops_buf2out_autovec_read_0_restart;
assign t_read[0] = output_sched_gen_0_valid_output;
assign loops_buf2out_autovec_read_1_step = t_read[1];
assign loops_sram2tb_mux_sel[1] = loops_buf2out_autovec_read_1_mux_sel_out;
assign loops_sram2tb_restart[1] = loops_buf2out_autovec_read_1_restart;
assign t_read[1] = output_sched_gen_1_valid_output;
for_loop_6_16 #(
  .CONFIG_WIDTH(5'h10),
  .ITERATOR_SUPPORT(4'h6))
loops_buf2out_autovec_read_0 (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_buf2out_autovec_read_0_dimensionality),
  .flush(flush),
  .ranges(loops_buf2out_autovec_read_0_ranges),
  .rst_n(rst_n),
  .step(loops_buf2out_autovec_read_0_step),
  .mux_sel_out(loops_buf2out_autovec_read_0_mux_sel_out),
  .restart(loops_buf2out_autovec_read_0_restart)
);

sched_gen_6_16 output_sched_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(output_sched_gen_0_enable),
  .finished(loops_buf2out_autovec_read_0_restart),
  .flush(flush),
  .mux_sel(loops_buf2out_autovec_read_0_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(output_sched_gen_0_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides(output_sched_gen_0_sched_addr_gen_strides),
  .valid_output(output_sched_gen_0_valid_output)
);

for_loop_6_16 #(
  .CONFIG_WIDTH(5'h10),
  .ITERATOR_SUPPORT(4'h6))
loops_buf2out_autovec_read_1 (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_buf2out_autovec_read_1_dimensionality),
  .flush(flush),
  .ranges(loops_buf2out_autovec_read_1_ranges),
  .rst_n(rst_n),
  .step(loops_buf2out_autovec_read_1_step),
  .mux_sel_out(loops_buf2out_autovec_read_1_mux_sel_out),
  .restart(loops_buf2out_autovec_read_1_restart)
);

sched_gen_6_16 output_sched_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(output_sched_gen_1_enable),
  .finished(loops_buf2out_autovec_read_1_restart),
  .flush(flush),
  .mux_sel(loops_buf2out_autovec_read_1_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(output_sched_gen_1_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides(output_sched_gen_1_sched_addr_gen_strides),
  .valid_output(output_sched_gen_1_valid_output)
);

endmodule   // strg_ub_sram_tb_shared

module strg_ub_tb_only (
  input logic clk,
  input logic clk_en,
  input logic [15:0] cycle_count,
  input logic flush,
  input logic [3:0] loops_buf2out_read_0_dimensionality,
  input logic [5:0] [15:0] loops_buf2out_read_0_ranges,
  input logic [3:0] loops_buf2out_read_1_dimensionality,
  input logic [5:0] [15:0] loops_buf2out_read_1_ranges,
  input logic [1:0] [2:0] loops_sram2tb_mux_sel,
  input logic [1:0] loops_sram2tb_restart,
  input logic rst_n,
  input logic [3:0] [15:0] sram_read_data,
  input logic [1:0] t_read,
  input logic [3:0] tb_read_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] tb_read_addr_gen_0_strides,
  input logic [3:0] tb_read_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] tb_read_addr_gen_1_strides,
  input logic tb_read_sched_gen_0_enable,
  input logic [15:0] tb_read_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] tb_read_sched_gen_0_sched_addr_gen_strides,
  input logic tb_read_sched_gen_1_enable,
  input logic [15:0] tb_read_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] tb_read_sched_gen_1_sched_addr_gen_strides,
  input logic [3:0] tb_write_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] tb_write_addr_gen_0_strides,
  input logic [3:0] tb_write_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] tb_write_addr_gen_1_strides,
  output logic [1:0] accessor_output,
  output logic [1:0] [15:0] data_out
);

logic [2:0] loops_buf2out_read_0_mux_sel_out;
logic loops_buf2out_read_0_restart;
logic loops_buf2out_read_0_step;
logic [2:0] loops_buf2out_read_1_mux_sel_out;
logic loops_buf2out_read_1_restart;
logic loops_buf2out_read_1_step;
logic [1:0][2:0] mux_sel_d1;
logic [1:0] restart_d1;
logic [1:0] t_read_d1;
logic [1:0][1:0][3:0][15:0] tb;
logic [1:0] tb_read;
logic [1:0][2:0] tb_read_addr;
logic [3:0] tb_read_addr_gen_0_addr_out;
logic tb_read_addr_gen_0_step;
logic [3:0] tb_read_addr_gen_1_addr_out;
logic tb_read_addr_gen_1_step;
logic tb_read_sched_gen_0_valid_output;
logic tb_read_sched_gen_1_valid_output;
logic [1:0][2:0] tb_write_addr;
logic [3:0] tb_write_addr_gen_0_addr_out;
logic [2:0] tb_write_addr_gen_0_mux_sel;
logic tb_write_addr_gen_0_restart;
logic tb_write_addr_gen_0_step;
logic [3:0] tb_write_addr_gen_1_addr_out;
logic [2:0] tb_write_addr_gen_1_mux_sel;
logic tb_write_addr_gen_1_restart;
logic tb_write_addr_gen_1_step;
assign accessor_output = tb_read;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    t_read_d1[0] <= 1'h0;
    mux_sel_d1[0] <= 3'h0;
    restart_d1[0] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      t_read_d1[0] <= 1'h0;
      mux_sel_d1[0] <= 3'h0;
      restart_d1[0] <= 1'h0;
    end
    else begin
      t_read_d1[0] <= t_read[0];
      mux_sel_d1[0] <= loops_sram2tb_mux_sel[0];
      restart_d1[0] <= loops_sram2tb_restart[0];
    end
  end
end

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    t_read_d1[1] <= 1'h0;
    mux_sel_d1[1] <= 3'h0;
    restart_d1[1] <= 1'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      t_read_d1[1] <= 1'h0;
      mux_sel_d1[1] <= 3'h0;
      restart_d1[1] <= 1'h0;
    end
    else begin
      t_read_d1[1] <= t_read[1];
      mux_sel_d1[1] <= loops_sram2tb_mux_sel[1];
      restart_d1[1] <= loops_sram2tb_restart[1];
    end
  end
end
assign tb_write_addr_gen_0_step = t_read_d1[0];
assign tb_write_addr_gen_0_mux_sel = mux_sel_d1[0];
assign tb_write_addr_gen_0_restart = restart_d1[0];
assign tb_write_addr[0] = tb_write_addr_gen_0_addr_out[2:0];

always_ff @(posedge clk) begin
  if (clk_en) begin
    if (t_read_d1[0]) begin
      tb[0][tb_write_addr[0][0]] <= sram_read_data;
    end
  end
end
assign loops_buf2out_read_0_step = tb_read[0];
assign tb_read_addr_gen_0_step = tb_read[0];
assign tb_read_addr[0] = tb_read_addr_gen_0_addr_out[2:0];
assign tb_read[0] = tb_read_sched_gen_0_valid_output;
always_comb begin
  data_out[0] = tb[0][tb_read_addr[0][2]][tb_read_addr[0][1:0]];
end
assign tb_write_addr_gen_1_step = t_read_d1[1];
assign tb_write_addr_gen_1_mux_sel = mux_sel_d1[1];
assign tb_write_addr_gen_1_restart = restart_d1[1];
assign tb_write_addr[1] = tb_write_addr_gen_1_addr_out[2:0];

always_ff @(posedge clk) begin
  if (clk_en) begin
    if (t_read_d1[1]) begin
      tb[1][tb_write_addr[1][0]] <= sram_read_data;
    end
  end
end
assign loops_buf2out_read_1_step = tb_read[1];
assign tb_read_addr_gen_1_step = tb_read[1];
assign tb_read_addr[1] = tb_read_addr_gen_1_addr_out[2:0];
assign tb_read[1] = tb_read_sched_gen_1_valid_output;
always_comb begin
  data_out[1] = tb[1][tb_read_addr[1][2]][tb_read_addr[1][1:0]];
end
addr_gen_6_4 tb_write_addr_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(tb_write_addr_gen_0_mux_sel),
  .restart(tb_write_addr_gen_0_restart),
  .rst_n(rst_n),
  .starting_addr(tb_write_addr_gen_0_starting_addr),
  .step(tb_write_addr_gen_0_step),
  .strides(tb_write_addr_gen_0_strides),
  .addr_out(tb_write_addr_gen_0_addr_out)
);

for_loop_6_16 #(
  .CONFIG_WIDTH(5'h10),
  .ITERATOR_SUPPORT(4'h6))
loops_buf2out_read_0 (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_buf2out_read_0_dimensionality),
  .flush(flush),
  .ranges(loops_buf2out_read_0_ranges),
  .rst_n(rst_n),
  .step(loops_buf2out_read_0_step),
  .mux_sel_out(loops_buf2out_read_0_mux_sel_out),
  .restart(loops_buf2out_read_0_restart)
);

addr_gen_6_4 tb_read_addr_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(loops_buf2out_read_0_mux_sel_out),
  .restart(loops_buf2out_read_0_restart),
  .rst_n(rst_n),
  .starting_addr(tb_read_addr_gen_0_starting_addr),
  .step(tb_read_addr_gen_0_step),
  .strides(tb_read_addr_gen_0_strides),
  .addr_out(tb_read_addr_gen_0_addr_out)
);

sched_gen_6_16 tb_read_sched_gen_0 (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(tb_read_sched_gen_0_enable),
  .finished(loops_buf2out_read_0_restart),
  .flush(flush),
  .mux_sel(loops_buf2out_read_0_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(tb_read_sched_gen_0_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides(tb_read_sched_gen_0_sched_addr_gen_strides),
  .valid_output(tb_read_sched_gen_0_valid_output)
);

addr_gen_6_4 tb_write_addr_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(tb_write_addr_gen_1_mux_sel),
  .restart(tb_write_addr_gen_1_restart),
  .rst_n(rst_n),
  .starting_addr(tb_write_addr_gen_1_starting_addr),
  .step(tb_write_addr_gen_1_step),
  .strides(tb_write_addr_gen_1_strides),
  .addr_out(tb_write_addr_gen_1_addr_out)
);

for_loop_6_16 #(
  .CONFIG_WIDTH(5'h10),
  .ITERATOR_SUPPORT(4'h6))
loops_buf2out_read_1 (
  .clk(clk),
  .clk_en(clk_en),
  .dimensionality(loops_buf2out_read_1_dimensionality),
  .flush(flush),
  .ranges(loops_buf2out_read_1_ranges),
  .rst_n(rst_n),
  .step(loops_buf2out_read_1_step),
  .mux_sel_out(loops_buf2out_read_1_mux_sel_out),
  .restart(loops_buf2out_read_1_restart)
);

addr_gen_6_4 tb_read_addr_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .flush(flush),
  .mux_sel(loops_buf2out_read_1_mux_sel_out),
  .restart(loops_buf2out_read_1_restart),
  .rst_n(rst_n),
  .starting_addr(tb_read_addr_gen_1_starting_addr),
  .step(tb_read_addr_gen_1_step),
  .strides(tb_read_addr_gen_1_strides),
  .addr_out(tb_read_addr_gen_1_addr_out)
);

sched_gen_6_16 tb_read_sched_gen_1 (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .enable(tb_read_sched_gen_1_enable),
  .finished(loops_buf2out_read_1_restart),
  .flush(flush),
  .mux_sel(loops_buf2out_read_1_mux_sel_out),
  .rst_n(rst_n),
  .sched_addr_gen_starting_addr(tb_read_sched_gen_1_sched_addr_gen_starting_addr),
  .sched_addr_gen_strides(tb_read_sched_gen_1_sched_addr_gen_strides),
  .valid_output(tb_read_sched_gen_1_valid_output)
);

endmodule   // strg_ub_tb_only

module strg_ub_vec (
  input logic [3:0] agg_only_agg_read_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] agg_only_agg_read_addr_gen_0_strides,
  input logic [3:0] agg_only_agg_read_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] agg_only_agg_read_addr_gen_1_strides,
  input logic [3:0] agg_only_agg_write_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] agg_only_agg_write_addr_gen_0_strides,
  input logic [3:0] agg_only_agg_write_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] agg_only_agg_write_addr_gen_1_strides,
  input logic agg_only_agg_write_sched_gen_0_enable,
  input logic [15:0] agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] agg_only_agg_write_sched_gen_0_sched_addr_gen_strides,
  input logic agg_only_agg_write_sched_gen_1_enable,
  input logic [15:0] agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] agg_only_agg_write_sched_gen_1_sched_addr_gen_strides,
  input logic [3:0] agg_only_loops_in2buf_0_dimensionality,
  input logic [5:0] [15:0] agg_only_loops_in2buf_0_ranges,
  input logic [3:0] agg_only_loops_in2buf_1_dimensionality,
  input logic [5:0] [15:0] agg_only_loops_in2buf_1_ranges,
  input logic agg_sram_shared_agg_read_sched_gen_0_enable,
  input logic [15:0] agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides,
  input logic agg_sram_shared_agg_read_sched_gen_1_enable,
  input logic [15:0] agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides,
  input logic [3:0] agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality,
  input logic [5:0] [15:0] agg_sram_shared_loops_in2buf_autovec_write_0_ranges,
  input logic [3:0] agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality,
  input logic [5:0] [15:0] agg_sram_shared_loops_in2buf_autovec_write_1_ranges,
  input logic clk,
  input logic clk_en,
  input logic [3:0] [15:0] data_from_strg,
  input logic [1:0] [15:0] data_in,
  input logic flush,
  input logic rst_n,
  input logic [8:0] sram_only_input_addr_gen_0_starting_addr,
  input logic [5:0] [8:0] sram_only_input_addr_gen_0_strides,
  input logic [8:0] sram_only_input_addr_gen_1_starting_addr,
  input logic [5:0] [8:0] sram_only_input_addr_gen_1_strides,
  input logic [8:0] sram_only_output_addr_gen_0_starting_addr,
  input logic [5:0] [8:0] sram_only_output_addr_gen_0_strides,
  input logic [8:0] sram_only_output_addr_gen_1_starting_addr,
  input logic [5:0] [8:0] sram_only_output_addr_gen_1_strides,
  input logic [3:0] sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality,
  input logic [5:0] [15:0] sram_tb_shared_loops_buf2out_autovec_read_0_ranges,
  input logic [3:0] sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality,
  input logic [5:0] [15:0] sram_tb_shared_loops_buf2out_autovec_read_1_ranges,
  input logic sram_tb_shared_output_sched_gen_0_enable,
  input logic [15:0] sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides,
  input logic sram_tb_shared_output_sched_gen_1_enable,
  input logic [15:0] sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides,
  input logic [3:0] tb_only_loops_buf2out_read_0_dimensionality,
  input logic [5:0] [15:0] tb_only_loops_buf2out_read_0_ranges,
  input logic [3:0] tb_only_loops_buf2out_read_1_dimensionality,
  input logic [5:0] [15:0] tb_only_loops_buf2out_read_1_ranges,
  input logic [3:0] tb_only_tb_read_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] tb_only_tb_read_addr_gen_0_strides,
  input logic [3:0] tb_only_tb_read_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] tb_only_tb_read_addr_gen_1_strides,
  input logic tb_only_tb_read_sched_gen_0_enable,
  input logic [15:0] tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] tb_only_tb_read_sched_gen_0_sched_addr_gen_strides,
  input logic tb_only_tb_read_sched_gen_1_enable,
  input logic [15:0] tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr,
  input logic [5:0] [15:0] tb_only_tb_read_sched_gen_1_sched_addr_gen_strides,
  input logic [3:0] tb_only_tb_write_addr_gen_0_starting_addr,
  input logic [5:0] [3:0] tb_only_tb_write_addr_gen_0_strides,
  input logic [3:0] tb_only_tb_write_addr_gen_1_starting_addr,
  input logic [5:0] [3:0] tb_only_tb_write_addr_gen_1_strides,
  output logic [1:0] accessor_output,
  output logic [8:0] addr_out,
  output logic cen_to_strg,
  output logic [1:0] [15:0] data_out,
  output logic [3:0] [15:0] data_to_strg,
  output logic wen_to_strg
);

logic [1:0][3:0][15:0] agg_only_agg_data_out;
logic [1:0] agg_only_agg_read;
logic [1:0][2:0] agg_only_floop_mux_sel;
logic [1:0] agg_only_floop_restart;
logic [1:0] agg_sram_shared_agg_read_out;
logic [1:0][2:0] agg_sram_shared_floop_mux_sel;
logic [1:0] agg_sram_shared_floop_restart;
logic [15:0] cycle_count;
logic [1:0][2:0] sram_only_loops_sram2tb_mux_sel;
logic [1:0] sram_only_loops_sram2tb_restart;
logic [1:0] sram_only_t_read;
logic [1:0][2:0] sram_tb_shared_loops_sram2tb_mux_sel;
logic [1:0] sram_tb_shared_loops_sram2tb_restart;
logic [1:0] sram_tb_shared_t_read_out;

always_ff @(posedge clk, negedge rst_n) begin
  if (~rst_n) begin
    cycle_count <= 16'h0;
  end
  else if (clk_en) begin
    if (flush) begin
      cycle_count <= 16'h0;
    end
    else if (1'h1) begin
      cycle_count <= cycle_count + 16'h1;
    end
  end
end
assign agg_only_agg_read = agg_sram_shared_agg_read_out;
assign agg_only_floop_mux_sel = agg_sram_shared_floop_mux_sel;
assign agg_only_floop_restart = agg_sram_shared_floop_restart;
assign sram_only_loops_sram2tb_mux_sel = sram_tb_shared_loops_sram2tb_mux_sel;
assign sram_only_loops_sram2tb_restart = sram_tb_shared_loops_sram2tb_restart;
assign sram_only_t_read = sram_tb_shared_t_read_out;
strg_ub_agg_only agg_only (
  .agg_read(agg_only_agg_read),
  .agg_read_addr_gen_0_starting_addr(agg_only_agg_read_addr_gen_0_starting_addr),
  .agg_read_addr_gen_0_strides(agg_only_agg_read_addr_gen_0_strides),
  .agg_read_addr_gen_1_starting_addr(agg_only_agg_read_addr_gen_1_starting_addr),
  .agg_read_addr_gen_1_strides(agg_only_agg_read_addr_gen_1_strides),
  .agg_write_addr_gen_0_starting_addr(agg_only_agg_write_addr_gen_0_starting_addr),
  .agg_write_addr_gen_0_strides(agg_only_agg_write_addr_gen_0_strides),
  .agg_write_addr_gen_1_starting_addr(agg_only_agg_write_addr_gen_1_starting_addr),
  .agg_write_addr_gen_1_strides(agg_only_agg_write_addr_gen_1_strides),
  .agg_write_sched_gen_0_enable(agg_only_agg_write_sched_gen_0_enable),
  .agg_write_sched_gen_0_sched_addr_gen_starting_addr(agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr),
  .agg_write_sched_gen_0_sched_addr_gen_strides(agg_only_agg_write_sched_gen_0_sched_addr_gen_strides),
  .agg_write_sched_gen_1_enable(agg_only_agg_write_sched_gen_1_enable),
  .agg_write_sched_gen_1_sched_addr_gen_starting_addr(agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr),
  .agg_write_sched_gen_1_sched_addr_gen_strides(agg_only_agg_write_sched_gen_1_sched_addr_gen_strides),
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .data_in(data_in),
  .floop_mux_sel(agg_only_floop_mux_sel),
  .floop_restart(agg_only_floop_restart),
  .flush(flush),
  .loops_in2buf_0_dimensionality(agg_only_loops_in2buf_0_dimensionality),
  .loops_in2buf_0_ranges(agg_only_loops_in2buf_0_ranges),
  .loops_in2buf_1_dimensionality(agg_only_loops_in2buf_1_dimensionality),
  .loops_in2buf_1_ranges(agg_only_loops_in2buf_1_ranges),
  .rst_n(rst_n),
  .agg_data_out(agg_only_agg_data_out)
);

strg_ub_agg_sram_shared agg_sram_shared (
  .agg_read_sched_gen_0_enable(agg_sram_shared_agg_read_sched_gen_0_enable),
  .agg_read_sched_gen_0_sched_addr_gen_starting_addr(agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr),
  .agg_read_sched_gen_0_sched_addr_gen_strides(agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides),
  .agg_read_sched_gen_1_enable(agg_sram_shared_agg_read_sched_gen_1_enable),
  .agg_read_sched_gen_1_sched_addr_gen_starting_addr(agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr),
  .agg_read_sched_gen_1_sched_addr_gen_strides(agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides),
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .flush(flush),
  .loops_in2buf_autovec_write_0_dimensionality(agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality),
  .loops_in2buf_autovec_write_0_ranges(agg_sram_shared_loops_in2buf_autovec_write_0_ranges),
  .loops_in2buf_autovec_write_1_dimensionality(agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality),
  .loops_in2buf_autovec_write_1_ranges(agg_sram_shared_loops_in2buf_autovec_write_1_ranges),
  .rst_n(rst_n),
  .agg_read_out(agg_sram_shared_agg_read_out),
  .floop_mux_sel(agg_sram_shared_floop_mux_sel),
  .floop_restart(agg_sram_shared_floop_restart)
);

strg_ub_sram_only sram_only (
  .agg_data_out(agg_only_agg_data_out),
  .agg_read(agg_sram_shared_agg_read_out),
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .floop_mux_sel(agg_sram_shared_floop_mux_sel),
  .floop_restart(agg_sram_shared_floop_restart),
  .flush(flush),
  .input_addr_gen_0_starting_addr(sram_only_input_addr_gen_0_starting_addr),
  .input_addr_gen_0_strides(sram_only_input_addr_gen_0_strides),
  .input_addr_gen_1_starting_addr(sram_only_input_addr_gen_1_starting_addr),
  .input_addr_gen_1_strides(sram_only_input_addr_gen_1_strides),
  .loops_sram2tb_mux_sel(sram_only_loops_sram2tb_mux_sel),
  .loops_sram2tb_restart(sram_only_loops_sram2tb_restart),
  .output_addr_gen_0_starting_addr(sram_only_output_addr_gen_0_starting_addr),
  .output_addr_gen_0_strides(sram_only_output_addr_gen_0_strides),
  .output_addr_gen_1_starting_addr(sram_only_output_addr_gen_1_starting_addr),
  .output_addr_gen_1_strides(sram_only_output_addr_gen_1_strides),
  .rst_n(rst_n),
  .t_read(sram_only_t_read),
  .addr_to_sram(addr_out),
  .cen_to_sram(cen_to_strg),
  .data_to_sram(data_to_strg),
  .wen_to_sram(wen_to_strg)
);

strg_ub_sram_tb_shared sram_tb_shared (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .flush(flush),
  .loops_buf2out_autovec_read_0_dimensionality(sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality),
  .loops_buf2out_autovec_read_0_ranges(sram_tb_shared_loops_buf2out_autovec_read_0_ranges),
  .loops_buf2out_autovec_read_1_dimensionality(sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality),
  .loops_buf2out_autovec_read_1_ranges(sram_tb_shared_loops_buf2out_autovec_read_1_ranges),
  .output_sched_gen_0_enable(sram_tb_shared_output_sched_gen_0_enable),
  .output_sched_gen_0_sched_addr_gen_starting_addr(sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr),
  .output_sched_gen_0_sched_addr_gen_strides(sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides),
  .output_sched_gen_1_enable(sram_tb_shared_output_sched_gen_1_enable),
  .output_sched_gen_1_sched_addr_gen_starting_addr(sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr),
  .output_sched_gen_1_sched_addr_gen_strides(sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides),
  .rst_n(rst_n),
  .loops_sram2tb_mux_sel(sram_tb_shared_loops_sram2tb_mux_sel),
  .loops_sram2tb_restart(sram_tb_shared_loops_sram2tb_restart),
  .t_read_out(sram_tb_shared_t_read_out)
);

strg_ub_tb_only tb_only (
  .clk(clk),
  .clk_en(clk_en),
  .cycle_count(cycle_count),
  .flush(flush),
  .loops_buf2out_read_0_dimensionality(tb_only_loops_buf2out_read_0_dimensionality),
  .loops_buf2out_read_0_ranges(tb_only_loops_buf2out_read_0_ranges),
  .loops_buf2out_read_1_dimensionality(tb_only_loops_buf2out_read_1_dimensionality),
  .loops_buf2out_read_1_ranges(tb_only_loops_buf2out_read_1_ranges),
  .loops_sram2tb_mux_sel(sram_tb_shared_loops_sram2tb_mux_sel),
  .loops_sram2tb_restart(sram_tb_shared_loops_sram2tb_restart),
  .rst_n(rst_n),
  .sram_read_data(data_from_strg),
  .t_read(sram_tb_shared_t_read_out),
  .tb_read_addr_gen_0_starting_addr(tb_only_tb_read_addr_gen_0_starting_addr),
  .tb_read_addr_gen_0_strides(tb_only_tb_read_addr_gen_0_strides),
  .tb_read_addr_gen_1_starting_addr(tb_only_tb_read_addr_gen_1_starting_addr),
  .tb_read_addr_gen_1_strides(tb_only_tb_read_addr_gen_1_strides),
  .tb_read_sched_gen_0_enable(tb_only_tb_read_sched_gen_0_enable),
  .tb_read_sched_gen_0_sched_addr_gen_starting_addr(tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr),
  .tb_read_sched_gen_0_sched_addr_gen_strides(tb_only_tb_read_sched_gen_0_sched_addr_gen_strides),
  .tb_read_sched_gen_1_enable(tb_only_tb_read_sched_gen_1_enable),
  .tb_read_sched_gen_1_sched_addr_gen_starting_addr(tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr),
  .tb_read_sched_gen_1_sched_addr_gen_strides(tb_only_tb_read_sched_gen_1_sched_addr_gen_strides),
  .tb_write_addr_gen_0_starting_addr(tb_only_tb_write_addr_gen_0_starting_addr),
  .tb_write_addr_gen_0_strides(tb_only_tb_write_addr_gen_0_strides),
  .tb_write_addr_gen_1_starting_addr(tb_only_tb_write_addr_gen_1_starting_addr),
  .tb_write_addr_gen_1_strides(tb_only_tb_write_addr_gen_1_strides),
  .accessor_output(accessor_output),
  .data_out(data_out)
);

endmodule   // strg_ub_vec


module LUT (
    input [7:0] lut,
    input bit0,
    input bit1,
    input bit2,
    output O,
    input CLK,
    input ASYNCRESET
);
wire bit_const_0_None_out;
wire [7:0] const_1_8_out;
wire [7:0] magma_Bits_8_and_inst0_out;
wire [7:0] magma_Bits_8_lshr_inst0_out;
corebit_const #(
    .value(1'b0)
) bit_const_0_None (
    .out(bit_const_0_None_out)
);
coreir_const #(
    .value(8'h01),
    .width(8)
) const_1_8 (
    .out(const_1_8_out)
);
coreir_and #(
    .width(8)
) magma_Bits_8_and_inst0 (
    .in0(magma_Bits_8_lshr_inst0_out),
    .in1(const_1_8_out),
    .out(magma_Bits_8_and_inst0_out)
);
wire [7:0] magma_Bits_8_lshr_inst0_in1;
assign magma_Bits_8_lshr_inst0_in1 = {bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit_const_0_None_out,bit2,bit1,bit0};
coreir_lshr #(
    .width(8)
) magma_Bits_8_lshr_inst0 (
    .in0(lut),
    .in1(magma_Bits_8_lshr_inst0_in1),
    .out(magma_Bits_8_lshr_inst0_out)
);
assign O = magma_Bits_8_and_inst0_out[0];
endmodule

module LTE (
    input [0:0] signed_,
    input [15:0] a,
    input [15:0] b,
    output [15:0] O0,
    output O1,
    output O2,
    output O3,
    output O4,
    output O5,
    input CLK,
    input ASYNCRESET
);
wire [0:0] Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [15:0] Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire bit_const_0_None_out;
wire [15:0] const_0_16_out;
wire [0:0] const_1_1_out;
wire magma_Bits_16_eq_inst0_out;
wire magma_Bits_16_sle_inst0_out;
wire magma_Bits_16_ule_inst0_out;
wire magma_Bits_1_eq_inst0_out;
coreir_mux #(
    .width(1)
) Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(magma_Bits_16_ule_inst0_out),
    .in1(magma_Bits_16_sle_inst0_out),
    .sel(magma_Bits_1_eq_inst0_out),
    .out(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(b),
    .in1(a),
    .sel(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .out(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
corebit_const #(
    .value(1'b0)
) bit_const_0_None (
    .out(bit_const_0_None_out)
);
coreir_const #(
    .value(16'h0000),
    .width(16)
) const_0_16 (
    .out(const_0_16_out)
);
coreir_const #(
    .value(1'h1),
    .width(1)
) const_1_1 (
    .out(const_1_1_out)
);
coreir_eq #(
    .width(16)
) magma_Bits_16_eq_inst0 (
    .in0(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(const_0_16_out),
    .out(magma_Bits_16_eq_inst0_out)
);
coreir_sle #(
    .width(16)
) magma_Bits_16_sle_inst0 (
    .in0(a),
    .in1(b),
    .out(magma_Bits_16_sle_inst0_out)
);
coreir_ule #(
    .width(16)
) magma_Bits_16_ule_inst0 (
    .in0(a),
    .in1(b),
    .out(magma_Bits_16_ule_inst0_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst0 (
    .in0(signed_),
    .in1(const_1_1_out),
    .out(magma_Bits_1_eq_inst0_out)
);
assign O0 = Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign O1 = Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign O2 = magma_Bits_16_eq_inst0_out;
assign O3 = Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out[15];
assign O4 = bit_const_0_None_out;
assign O5 = bit_const_0_None_out;
endmodule

module GTE (
    input [0:0] signed_,
    input [15:0] a,
    input [15:0] b,
    output [15:0] O0,
    output O1,
    output O2,
    output O3,
    output O4,
    output O5,
    input CLK,
    input ASYNCRESET
);
wire [0:0] Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [15:0] Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire bit_const_0_None_out;
wire [15:0] const_0_16_out;
wire [0:0] const_1_1_out;
wire magma_Bits_16_eq_inst0_out;
wire magma_Bits_16_sge_inst0_out;
wire magma_Bits_16_uge_inst0_out;
wire magma_Bits_1_eq_inst0_out;
coreir_mux #(
    .width(1)
) Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(magma_Bits_16_uge_inst0_out),
    .in1(magma_Bits_16_sge_inst0_out),
    .sel(magma_Bits_1_eq_inst0_out),
    .out(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(b),
    .in1(a),
    .sel(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .out(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
corebit_const #(
    .value(1'b0)
) bit_const_0_None (
    .out(bit_const_0_None_out)
);
coreir_const #(
    .value(16'h0000),
    .width(16)
) const_0_16 (
    .out(const_0_16_out)
);
coreir_const #(
    .value(1'h1),
    .width(1)
) const_1_1 (
    .out(const_1_1_out)
);
coreir_eq #(
    .width(16)
) magma_Bits_16_eq_inst0 (
    .in0(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(const_0_16_out),
    .out(magma_Bits_16_eq_inst0_out)
);
coreir_sge #(
    .width(16)
) magma_Bits_16_sge_inst0 (
    .in0(a),
    .in1(b),
    .out(magma_Bits_16_sge_inst0_out)
);
coreir_uge #(
    .width(16)
) magma_Bits_16_uge_inst0 (
    .in0(a),
    .in1(b),
    .out(magma_Bits_16_uge_inst0_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst0 (
    .in0(signed_),
    .in1(const_1_1_out),
    .out(magma_Bits_1_eq_inst0_out)
);
assign O0 = Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign O1 = Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign O2 = magma_Bits_16_eq_inst0_out;
assign O3 = Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out[15];
assign O4 = bit_const_0_None_out;
assign O5 = bit_const_0_None_out;
endmodule

module Decode98 (
    input [7:0] I,
    output O
);
wire [7:0] const_9_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h09),
    .width(8)
) const_9_8 (
    .out(const_9_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_9_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode88 (
    input [7:0] I,
    output O
);
wire [7:0] const_8_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h08),
    .width(8)
) const_8_8 (
    .out(const_8_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_8_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode78 (
    input [7:0] I,
    output O
);
wire [7:0] const_7_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h07),
    .width(8)
) const_7_8 (
    .out(const_7_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_7_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode68 (
    input [7:0] I,
    output O
);
wire [7:0] const_6_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h06),
    .width(8)
) const_6_8 (
    .out(const_6_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_6_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode58 (
    input [7:0] I,
    output O
);
wire [7:0] const_5_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h05),
    .width(8)
) const_5_8 (
    .out(const_5_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_5_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode48 (
    input [7:0] I,
    output O
);
wire [7:0] const_4_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h04),
    .width(8)
) const_4_8 (
    .out(const_4_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_4_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode38 (
    input [7:0] I,
    output O
);
wire [7:0] const_3_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h03),
    .width(8)
) const_3_8 (
    .out(const_3_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_3_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode28 (
    input [7:0] I,
    output O
);
wire [7:0] const_2_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h02),
    .width(8)
) const_2_8 (
    .out(const_2_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_2_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode18 (
    input [7:0] I,
    output O
);
wire [7:0] const_1_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h01),
    .width(8)
) const_1_8 (
    .out(const_1_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_1_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode158 (
    input [7:0] I,
    output O
);
wire [7:0] const_15_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h0f),
    .width(8)
) const_15_8 (
    .out(const_15_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_15_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode148 (
    input [7:0] I,
    output O
);
wire [7:0] const_14_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h0e),
    .width(8)
) const_14_8 (
    .out(const_14_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_14_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode138 (
    input [7:0] I,
    output O
);
wire [7:0] const_13_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h0d),
    .width(8)
) const_13_8 (
    .out(const_13_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_13_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode128 (
    input [7:0] I,
    output O
);
wire [7:0] const_12_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h0c),
    .width(8)
) const_12_8 (
    .out(const_12_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_12_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode118 (
    input [7:0] I,
    output O
);
wire [7:0] const_11_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h0b),
    .width(8)
) const_11_8 (
    .out(const_11_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_11_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode108 (
    input [7:0] I,
    output O
);
wire [7:0] const_10_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h0a),
    .width(8)
) const_10_8 (
    .out(const_10_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_10_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module Decode08 (
    input [7:0] I,
    output O
);
wire [7:0] const_0_8_out;
wire coreir_eq_8_inst0_out;
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
coreir_eq #(
    .width(8)
) coreir_eq_8_inst0 (
    .in0(I),
    .in1(const_0_8_out),
    .out(coreir_eq_8_inst0_out)
);
assign O = coreir_eq_8_inst0_out;
endmodule

module ConfigRegister_5_8_32_0 (
    input clk,
    input reset,
    output [4:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [4:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_5_inst0_O;
wire [7:0] const_0_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_5 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_5_inst0 (
    .I(config_data[4:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_5_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_0_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_5_inst0_O;
endmodule

module ConfigRegister_4_8_32_3 (
    input clk,
    input reset,
    output [3:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [3:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_4_inst0_O;
wire [7:0] const_3_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_4 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_4_inst0 (
    .I(config_data[3:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_4_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h03),
    .width(8)
) const_3_8 (
    .out(const_3_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_3_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_4_inst0_O;
endmodule

module ConfigRegister_32_8_32_9 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_9_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h09),
    .width(8)
) const_9_8 (
    .out(const_9_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_9_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_82 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_82_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h52),
    .width(8)
) const_82_8 (
    .out(const_82_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_82_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_81 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_81_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h51),
    .width(8)
) const_81_8 (
    .out(const_81_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_81_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_80 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_80_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h50),
    .width(8)
) const_80_8 (
    .out(const_80_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_80_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_8 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_8_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h08),
    .width(8)
) const_8_8 (
    .out(const_8_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_8_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_79 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_79_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h4f),
    .width(8)
) const_79_8 (
    .out(const_79_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_79_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_77 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_77_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h4d),
    .width(8)
) const_77_8 (
    .out(const_77_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_77_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_76 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_76_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h4c),
    .width(8)
) const_76_8 (
    .out(const_76_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_76_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_75 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_75_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h4b),
    .width(8)
) const_75_8 (
    .out(const_75_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_75_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_73 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_73_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h49),
    .width(8)
) const_73_8 (
    .out(const_73_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_73_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_72 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_72_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h48),
    .width(8)
) const_72_8 (
    .out(const_72_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_72_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_71 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_71_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h47),
    .width(8)
) const_71_8 (
    .out(const_71_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_71_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_70 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_70_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h46),
    .width(8)
) const_70_8 (
    .out(const_70_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_70_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_7 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_7_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h07),
    .width(8)
) const_7_8 (
    .out(const_7_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_7_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_68 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_68_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h44),
    .width(8)
) const_68_8 (
    .out(const_68_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_68_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_67 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_67_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h43),
    .width(8)
) const_67_8 (
    .out(const_67_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_67_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_66 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_66_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h42),
    .width(8)
) const_66_8 (
    .out(const_66_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_66_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_64 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_64_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h40),
    .width(8)
) const_64_8 (
    .out(const_64_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_64_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_63 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_63_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h3f),
    .width(8)
) const_63_8 (
    .out(const_63_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_63_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_62 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_62_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h3e),
    .width(8)
) const_62_8 (
    .out(const_62_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_62_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_60 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_60_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h3c),
    .width(8)
) const_60_8 (
    .out(const_60_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_60_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_6 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_6_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h06),
    .width(8)
) const_6_8 (
    .out(const_6_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_6_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_59 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_59_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h3b),
    .width(8)
) const_59_8 (
    .out(const_59_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_59_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_58 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_58_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h3a),
    .width(8)
) const_58_8 (
    .out(const_58_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_58_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_56 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_56_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h38),
    .width(8)
) const_56_8 (
    .out(const_56_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_56_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_55 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_55_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h37),
    .width(8)
) const_55_8 (
    .out(const_55_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_55_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_53 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_53_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h35),
    .width(8)
) const_53_8 (
    .out(const_53_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_53_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_52 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_52_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h34),
    .width(8)
) const_52_8 (
    .out(const_52_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_52_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_51 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_51_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h33),
    .width(8)
) const_51_8 (
    .out(const_51_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_51_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_5 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_5_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h05),
    .width(8)
) const_5_8 (
    .out(const_5_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_5_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_40 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_40_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h28),
    .width(8)
) const_40_8 (
    .out(const_40_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_40_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_39 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_39_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h27),
    .width(8)
) const_39_8 (
    .out(const_39_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_39_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_37 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_37_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h25),
    .width(8)
) const_37_8 (
    .out(const_37_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_37_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_36 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_36_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h24),
    .width(8)
) const_36_8 (
    .out(const_36_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_36_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_35 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_35_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h23),
    .width(8)
) const_35_8 (
    .out(const_35_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_35_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_33 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_33_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h21),
    .width(8)
) const_33_8 (
    .out(const_33_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_33_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_32 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_32_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h20),
    .width(8)
) const_32_8 (
    .out(const_32_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_32_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_31 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_31_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h1f),
    .width(8)
) const_31_8 (
    .out(const_31_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_31_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_3 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_3_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h03),
    .width(8)
) const_3_8 (
    .out(const_3_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_3_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_29 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_29_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h1d),
    .width(8)
) const_29_8 (
    .out(const_29_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_29_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_28 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_28_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h1c),
    .width(8)
) const_28_8 (
    .out(const_28_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_28_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_27 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_27_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h1b),
    .width(8)
) const_27_8 (
    .out(const_27_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_27_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_25 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_25_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h19),
    .width(8)
) const_25_8 (
    .out(const_25_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_25_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_24 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_24_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h18),
    .width(8)
) const_24_8 (
    .out(const_24_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_24_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_22 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_22_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h16),
    .width(8)
) const_22_8 (
    .out(const_22_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_22_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_21 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_21_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h15),
    .width(8)
) const_21_8 (
    .out(const_21_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_21_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_20 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_20_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h14),
    .width(8)
) const_20_8 (
    .out(const_20_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_20_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_2 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_2_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h02),
    .width(8)
) const_2_8 (
    .out(const_2_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_2_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_18 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_18_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h12),
    .width(8)
) const_18_8 (
    .out(const_18_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_18_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_17 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_17_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h11),
    .width(8)
) const_17_8 (
    .out(const_17_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_17_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_16 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_16_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h10),
    .width(8)
) const_16_8 (
    .out(const_16_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_16_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_14 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_14_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h0e),
    .width(8)
) const_14_8 (
    .out(const_14_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_14_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_13 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_13_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h0d),
    .width(8)
) const_13_8 (
    .out(const_13_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_13_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_12 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_12_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h0c),
    .width(8)
) const_12_8 (
    .out(const_12_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_12_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_10 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_10_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h0a),
    .width(8)
) const_10_8 (
    .out(const_10_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_10_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_1 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_1_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h01),
    .width(8)
) const_1_8 (
    .out(const_1_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_1_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module ConfigRegister_32_8_32_0 (
    input clk,
    input reset,
    output [31:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [31:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
wire [7:0] const_0_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0 (
    .I(config_data),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_0_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_32_inst0_O;
endmodule

module SB_ID0_5TRACKS_B1_MemCore (
    input [0:0] SB_T0_EAST_SB_IN_B1,
    output [0:0] SB_T0_EAST_SB_OUT_B1,
    input [0:0] SB_T0_NORTH_SB_IN_B1,
    output [0:0] SB_T0_NORTH_SB_OUT_B1,
    input [0:0] SB_T0_SOUTH_SB_IN_B1,
    output [0:0] SB_T0_SOUTH_SB_OUT_B1,
    input [0:0] SB_T0_WEST_SB_IN_B1,
    output [0:0] SB_T0_WEST_SB_OUT_B1,
    input [0:0] SB_T1_EAST_SB_IN_B1,
    output [0:0] SB_T1_EAST_SB_OUT_B1,
    input [0:0] SB_T1_NORTH_SB_IN_B1,
    output [0:0] SB_T1_NORTH_SB_OUT_B1,
    input [0:0] SB_T1_SOUTH_SB_IN_B1,
    output [0:0] SB_T1_SOUTH_SB_OUT_B1,
    input [0:0] SB_T1_WEST_SB_IN_B1,
    output [0:0] SB_T1_WEST_SB_OUT_B1,
    input [0:0] SB_T2_EAST_SB_IN_B1,
    output [0:0] SB_T2_EAST_SB_OUT_B1,
    input [0:0] SB_T2_NORTH_SB_IN_B1,
    output [0:0] SB_T2_NORTH_SB_OUT_B1,
    input [0:0] SB_T2_SOUTH_SB_IN_B1,
    output [0:0] SB_T2_SOUTH_SB_OUT_B1,
    input [0:0] SB_T2_WEST_SB_IN_B1,
    output [0:0] SB_T2_WEST_SB_OUT_B1,
    input [0:0] SB_T3_EAST_SB_IN_B1,
    output [0:0] SB_T3_EAST_SB_OUT_B1,
    input [0:0] SB_T3_NORTH_SB_IN_B1,
    output [0:0] SB_T3_NORTH_SB_OUT_B1,
    input [0:0] SB_T3_SOUTH_SB_IN_B1,
    output [0:0] SB_T3_SOUTH_SB_OUT_B1,
    input [0:0] SB_T3_WEST_SB_IN_B1,
    output [0:0] SB_T3_WEST_SB_OUT_B1,
    input [0:0] SB_T4_EAST_SB_IN_B1,
    output [0:0] SB_T4_EAST_SB_OUT_B1,
    input [0:0] SB_T4_NORTH_SB_IN_B1,
    output [0:0] SB_T4_NORTH_SB_OUT_B1,
    input [0:0] SB_T4_SOUTH_SB_IN_B1,
    output [0:0] SB_T4_SOUTH_SB_OUT_B1,
    input [0:0] SB_T4_WEST_SB_IN_B1,
    output [0:0] SB_T4_WEST_SB_OUT_B1,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    input [0:0] empty,
    input [0:0] full,
    output [31:0] read_config_data,
    input reset,
    input [0:0] sram_ready_out,
    input [0:0] stall,
    input [0:0] stencil_valid,
    input [0:0] valid_out_0,
    input [0:0] valid_out_1
);
wire [0:0] Invert1_inst0_out;
wire [0:0] MUX_SB_T0_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out;
wire [0:0] MUX_SB_T0_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out;
wire [0:0] MUX_SB_T0_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out;
wire [0:0] MUX_SB_T0_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out;
wire [0:0] MUX_SB_T1_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out;
wire [0:0] MUX_SB_T1_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out;
wire [0:0] MUX_SB_T1_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out;
wire [0:0] MUX_SB_T1_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out;
wire [0:0] MUX_SB_T2_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out;
wire [0:0] MUX_SB_T2_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out;
wire [0:0] MUX_SB_T2_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out;
wire [0:0] MUX_SB_T2_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out;
wire [0:0] MUX_SB_T3_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out;
wire [0:0] MUX_SB_T3_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out;
wire [0:0] MUX_SB_T3_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out;
wire [0:0] MUX_SB_T3_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out;
wire [0:0] MUX_SB_T4_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out;
wire [0:0] MUX_SB_T4_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out;
wire [0:0] MUX_SB_T4_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out;
wire [0:0] MUX_SB_T4_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out;
wire [31:0] MuxWrapper_4_32_inst0$Mux4x32_inst0$coreir_commonlib_mux4x32_inst0_out;
wire [1:0] MuxWrapper_4_32_inst0_S_in;
wire [0:0] REG_T0_EAST_B1_O;
wire [0:0] REG_T0_NORTH_B1_O;
wire [0:0] REG_T0_SOUTH_B1_O;
wire [0:0] REG_T0_WEST_B1_O;
wire [0:0] REG_T1_EAST_B1_O;
wire [0:0] REG_T1_NORTH_B1_O;
wire [0:0] REG_T1_SOUTH_B1_O;
wire [0:0] REG_T1_WEST_B1_O;
wire [0:0] REG_T2_EAST_B1_O;
wire [0:0] REG_T2_NORTH_B1_O;
wire [0:0] REG_T2_SOUTH_B1_O;
wire [0:0] REG_T2_WEST_B1_O;
wire [0:0] REG_T3_EAST_B1_O;
wire [0:0] REG_T3_NORTH_B1_O;
wire [0:0] REG_T3_SOUTH_B1_O;
wire [0:0] REG_T3_WEST_B1_O;
wire [0:0] REG_T4_EAST_B1_O;
wire [0:0] REG_T4_NORTH_B1_O;
wire [0:0] REG_T4_SOUTH_B1_O;
wire [0:0] REG_T4_WEST_B1_O;
wire [0:0] RMUX_T0_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T0_EAST_B1_sel_inst0_O;
wire [0:0] RMUX_T0_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T0_NORTH_B1_sel_inst0_O;
wire [0:0] RMUX_T0_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T0_SOUTH_B1_sel_inst0_O;
wire [0:0] RMUX_T0_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T0_WEST_B1_sel_inst0_O;
wire [0:0] RMUX_T1_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T1_EAST_B1_sel_inst0_O;
wire [0:0] RMUX_T1_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T1_NORTH_B1_sel_inst0_O;
wire [0:0] RMUX_T1_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T1_SOUTH_B1_sel_inst0_O;
wire [0:0] RMUX_T1_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T1_WEST_B1_sel_inst0_O;
wire [0:0] RMUX_T2_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T2_EAST_B1_sel_inst0_O;
wire [0:0] RMUX_T2_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T2_NORTH_B1_sel_inst0_O;
wire [0:0] RMUX_T2_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T2_SOUTH_B1_sel_inst0_O;
wire [0:0] RMUX_T2_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T2_WEST_B1_sel_inst0_O;
wire [0:0] RMUX_T3_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T3_EAST_B1_sel_inst0_O;
wire [0:0] RMUX_T3_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T3_NORTH_B1_sel_inst0_O;
wire [0:0] RMUX_T3_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T3_SOUTH_B1_sel_inst0_O;
wire [0:0] RMUX_T3_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T3_WEST_B1_sel_inst0_O;
wire [0:0] RMUX_T4_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T4_EAST_B1_sel_inst0_O;
wire [0:0] RMUX_T4_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T4_NORTH_B1_sel_inst0_O;
wire [0:0] RMUX_T4_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T4_SOUTH_B1_sel_inst0_O;
wire [0:0] RMUX_T4_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T4_WEST_B1_sel_inst0_O;
wire [3:0] SB_T0_EAST_SB_OUT_B1_sel_inst0_O;
wire [3:0] SB_T0_NORTH_SB_OUT_B1_sel_inst0_O;
wire [3:0] SB_T0_SOUTH_SB_OUT_B1_sel_inst0_O;
wire [3:0] SB_T0_WEST_SB_OUT_B1_sel_inst0_O;
wire [3:0] SB_T1_EAST_SB_OUT_B1_sel_inst0_O;
wire [3:0] SB_T1_NORTH_SB_OUT_B1_sel_inst0_O;
wire [3:0] SB_T1_SOUTH_SB_OUT_B1_sel_inst0_O;
wire [3:0] SB_T1_WEST_SB_OUT_B1_sel_inst0_O;
wire [3:0] SB_T2_EAST_SB_OUT_B1_sel_inst0_O;
wire [3:0] SB_T2_NORTH_SB_OUT_B1_sel_inst0_O;
wire [3:0] SB_T2_SOUTH_SB_OUT_B1_sel_inst0_O;
wire [3:0] SB_T2_WEST_SB_OUT_B1_sel_inst0_O;
wire [3:0] SB_T3_EAST_SB_OUT_B1_sel_inst0_O;
wire [3:0] SB_T3_NORTH_SB_OUT_B1_sel_inst0_O;
wire [3:0] SB_T3_SOUTH_SB_OUT_B1_sel_inst0_O;
wire [3:0] SB_T3_WEST_SB_OUT_B1_sel_inst0_O;
wire [3:0] SB_T4_EAST_SB_OUT_B1_sel_inst0_O;
wire [3:0] SB_T4_NORTH_SB_OUT_B1_sel_inst0_O;
wire [3:0] SB_T4_SOUTH_SB_OUT_B1_sel_inst0_O;
wire [3:0] SB_T4_WEST_SB_OUT_B1_sel_inst0_O;
wire [0:0] WIRE_SB_T0_EAST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T0_NORTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T0_SOUTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T0_WEST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T1_EAST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T1_NORTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T1_SOUTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T1_WEST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T2_EAST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T2_NORTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T2_SOUTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T2_WEST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T3_EAST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T3_NORTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T3_SOUTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T3_WEST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T4_EAST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T4_NORTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T4_SOUTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T4_WEST_SB_IN_B1_O;
wire ZextWrapper_4_32_inst0$bit_const_0_None_out;
wire [3:0] ZextWrapper_4_32_inst0$self_I_out;
wire [31:0] ZextWrapper_4_32_inst0$self_O_in;
wire [0:0] and1_inst0_out;
wire [0:0] and1_inst1_out;
wire [0:0] and1_inst10_out;
wire [0:0] and1_inst11_out;
wire [0:0] and1_inst12_out;
wire [0:0] and1_inst13_out;
wire [0:0] and1_inst14_out;
wire [0:0] and1_inst15_out;
wire [0:0] and1_inst16_out;
wire [0:0] and1_inst17_out;
wire [0:0] and1_inst18_out;
wire [0:0] and1_inst19_out;
wire [0:0] and1_inst2_out;
wire [0:0] and1_inst3_out;
wire [0:0] and1_inst4_out;
wire [0:0] and1_inst5_out;
wire [0:0] and1_inst6_out;
wire [0:0] and1_inst7_out;
wire [0:0] and1_inst8_out;
wire [0:0] and1_inst9_out;
wire [31:0] config_reg_0_O;
wire [31:0] config_reg_1_O;
wire [31:0] config_reg_2_O;
wire [3:0] config_reg_3_O;
wire [0:0] const_1_1_out;
wire coreir_eq_1_inst0_out;
wire coreir_eq_1_inst1_out;
wire coreir_eq_1_inst10_out;
wire coreir_eq_1_inst11_out;
wire coreir_eq_1_inst12_out;
wire coreir_eq_1_inst13_out;
wire coreir_eq_1_inst14_out;
wire coreir_eq_1_inst15_out;
wire coreir_eq_1_inst16_out;
wire coreir_eq_1_inst17_out;
wire coreir_eq_1_inst18_out;
wire coreir_eq_1_inst19_out;
wire coreir_eq_1_inst2_out;
wire coreir_eq_1_inst3_out;
wire coreir_eq_1_inst4_out;
wire coreir_eq_1_inst5_out;
wire coreir_eq_1_inst6_out;
wire coreir_eq_1_inst7_out;
wire coreir_eq_1_inst8_out;
wire coreir_eq_1_inst9_out;
wire [7:0] self_config_config_addr_out;
coreir_not #(
    .width(1)
) Invert1_inst0 (
    .in(stall),
    .out(Invert1_inst0_out)
);
commonlib_muxn__N9__width1 MUX_SB_T0_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0 (
    .in_data_0(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .in_data_3(empty),
    .in_data_4(full),
    .in_data_5(sram_ready_out),
    .in_data_6(stencil_valid),
    .in_data_7(valid_out_0),
    .in_data_8(valid_out_1),
    .in_sel(SB_T0_EAST_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T0_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out)
);
commonlib_muxn__N9__width1 MUX_SB_T0_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0 (
    .in_data_0(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .in_data_3(empty),
    .in_data_4(full),
    .in_data_5(sram_ready_out),
    .in_data_6(stencil_valid),
    .in_data_7(valid_out_0),
    .in_data_8(valid_out_1),
    .in_sel(SB_T0_NORTH_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T0_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out)
);
commonlib_muxn__N9__width1 MUX_SB_T0_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0 (
    .in_data_0(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .in_data_3(empty),
    .in_data_4(full),
    .in_data_5(sram_ready_out),
    .in_data_6(stencil_valid),
    .in_data_7(valid_out_0),
    .in_data_8(valid_out_1),
    .in_sel(SB_T0_SOUTH_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T0_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out)
);
commonlib_muxn__N9__width1 MUX_SB_T0_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0 (
    .in_data_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .in_data_3(empty),
    .in_data_4(full),
    .in_data_5(sram_ready_out),
    .in_data_6(stencil_valid),
    .in_data_7(valid_out_0),
    .in_data_8(valid_out_1),
    .in_sel(SB_T0_WEST_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T0_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out)
);
commonlib_muxn__N9__width1 MUX_SB_T1_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0 (
    .in_data_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .in_data_3(empty),
    .in_data_4(full),
    .in_data_5(sram_ready_out),
    .in_data_6(stencil_valid),
    .in_data_7(valid_out_0),
    .in_data_8(valid_out_1),
    .in_sel(SB_T1_EAST_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T1_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out)
);
commonlib_muxn__N9__width1 MUX_SB_T1_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0 (
    .in_data_0(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .in_data_3(empty),
    .in_data_4(full),
    .in_data_5(sram_ready_out),
    .in_data_6(stencil_valid),
    .in_data_7(valid_out_0),
    .in_data_8(valid_out_1),
    .in_sel(SB_T1_NORTH_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T1_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out)
);
commonlib_muxn__N9__width1 MUX_SB_T1_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0 (
    .in_data_0(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .in_data_3(empty),
    .in_data_4(full),
    .in_data_5(sram_ready_out),
    .in_data_6(stencil_valid),
    .in_data_7(valid_out_0),
    .in_data_8(valid_out_1),
    .in_sel(SB_T1_SOUTH_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T1_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out)
);
commonlib_muxn__N9__width1 MUX_SB_T1_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0 (
    .in_data_0(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .in_data_3(empty),
    .in_data_4(full),
    .in_data_5(sram_ready_out),
    .in_data_6(stencil_valid),
    .in_data_7(valid_out_0),
    .in_data_8(valid_out_1),
    .in_sel(SB_T1_WEST_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T1_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out)
);
commonlib_muxn__N9__width1 MUX_SB_T2_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0 (
    .in_data_0(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .in_data_3(empty),
    .in_data_4(full),
    .in_data_5(sram_ready_out),
    .in_data_6(stencil_valid),
    .in_data_7(valid_out_0),
    .in_data_8(valid_out_1),
    .in_sel(SB_T2_EAST_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T2_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out)
);
commonlib_muxn__N9__width1 MUX_SB_T2_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0 (
    .in_data_0(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .in_data_3(empty),
    .in_data_4(full),
    .in_data_5(sram_ready_out),
    .in_data_6(stencil_valid),
    .in_data_7(valid_out_0),
    .in_data_8(valid_out_1),
    .in_sel(SB_T2_NORTH_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T2_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out)
);
commonlib_muxn__N9__width1 MUX_SB_T2_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0 (
    .in_data_0(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .in_data_3(empty),
    .in_data_4(full),
    .in_data_5(sram_ready_out),
    .in_data_6(stencil_valid),
    .in_data_7(valid_out_0),
    .in_data_8(valid_out_1),
    .in_sel(SB_T2_SOUTH_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T2_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out)
);
commonlib_muxn__N9__width1 MUX_SB_T2_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0 (
    .in_data_0(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .in_data_3(empty),
    .in_data_4(full),
    .in_data_5(sram_ready_out),
    .in_data_6(stencil_valid),
    .in_data_7(valid_out_0),
    .in_data_8(valid_out_1),
    .in_sel(SB_T2_WEST_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T2_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out)
);
commonlib_muxn__N9__width1 MUX_SB_T3_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0 (
    .in_data_0(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .in_data_3(empty),
    .in_data_4(full),
    .in_data_5(sram_ready_out),
    .in_data_6(stencil_valid),
    .in_data_7(valid_out_0),
    .in_data_8(valid_out_1),
    .in_sel(SB_T3_EAST_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T3_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out)
);
commonlib_muxn__N9__width1 MUX_SB_T3_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0 (
    .in_data_0(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .in_data_3(empty),
    .in_data_4(full),
    .in_data_5(sram_ready_out),
    .in_data_6(stencil_valid),
    .in_data_7(valid_out_0),
    .in_data_8(valid_out_1),
    .in_sel(SB_T3_NORTH_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T3_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out)
);
commonlib_muxn__N9__width1 MUX_SB_T3_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0 (
    .in_data_0(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .in_data_3(empty),
    .in_data_4(full),
    .in_data_5(sram_ready_out),
    .in_data_6(stencil_valid),
    .in_data_7(valid_out_0),
    .in_data_8(valid_out_1),
    .in_sel(SB_T3_SOUTH_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T3_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out)
);
commonlib_muxn__N9__width1 MUX_SB_T3_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0 (
    .in_data_0(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .in_data_3(empty),
    .in_data_4(full),
    .in_data_5(sram_ready_out),
    .in_data_6(stencil_valid),
    .in_data_7(valid_out_0),
    .in_data_8(valid_out_1),
    .in_sel(SB_T3_WEST_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T3_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out)
);
commonlib_muxn__N9__width1 MUX_SB_T4_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0 (
    .in_data_0(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .in_data_3(empty),
    .in_data_4(full),
    .in_data_5(sram_ready_out),
    .in_data_6(stencil_valid),
    .in_data_7(valid_out_0),
    .in_data_8(valid_out_1),
    .in_sel(SB_T4_EAST_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T4_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out)
);
commonlib_muxn__N9__width1 MUX_SB_T4_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0 (
    .in_data_0(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .in_data_3(empty),
    .in_data_4(full),
    .in_data_5(sram_ready_out),
    .in_data_6(stencil_valid),
    .in_data_7(valid_out_0),
    .in_data_8(valid_out_1),
    .in_sel(SB_T4_NORTH_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T4_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out)
);
commonlib_muxn__N9__width1 MUX_SB_T4_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0 (
    .in_data_0(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .in_data_3(empty),
    .in_data_4(full),
    .in_data_5(sram_ready_out),
    .in_data_6(stencil_valid),
    .in_data_7(valid_out_0),
    .in_data_8(valid_out_1),
    .in_sel(SB_T4_SOUTH_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T4_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out)
);
commonlib_muxn__N9__width1 MUX_SB_T4_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0 (
    .in_data_0(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .in_data_3(empty),
    .in_data_4(full),
    .in_data_5(sram_ready_out),
    .in_data_6(stencil_valid),
    .in_data_7(valid_out_0),
    .in_data_8(valid_out_1),
    .in_sel(SB_T4_WEST_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T4_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out)
);
commonlib_muxn__N4__width32 MuxWrapper_4_32_inst0$Mux4x32_inst0$coreir_commonlib_mux4x32_inst0 (
    .in_data_0(config_reg_0_O),
    .in_data_1(config_reg_1_O),
    .in_data_2(config_reg_2_O),
    .in_data_3(ZextWrapper_4_32_inst0$self_O_in),
    .in_sel(MuxWrapper_4_32_inst0_S_in),
    .out(MuxWrapper_4_32_inst0$Mux4x32_inst0$coreir_commonlib_mux4x32_inst0_out)
);
mantle_wire__typeBitIn2 MuxWrapper_4_32_inst0_S (
    .in(MuxWrapper_4_32_inst0_S_in),
    .out(self_config_config_addr_out[1:0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T0_EAST_B1 (
    .I(MUX_SB_T0_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .O(REG_T0_EAST_B1_O),
    .CLK(clk),
    .CE(and1_inst2_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T0_NORTH_B1 (
    .I(MUX_SB_T0_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .O(REG_T0_NORTH_B1_O),
    .CLK(clk),
    .CE(and1_inst0_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T0_SOUTH_B1 (
    .I(MUX_SB_T0_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .O(REG_T0_SOUTH_B1_O),
    .CLK(clk),
    .CE(and1_inst1_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T0_WEST_B1 (
    .I(MUX_SB_T0_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .O(REG_T0_WEST_B1_O),
    .CLK(clk),
    .CE(and1_inst3_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T1_EAST_B1 (
    .I(MUX_SB_T1_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .O(REG_T1_EAST_B1_O),
    .CLK(clk),
    .CE(and1_inst6_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T1_NORTH_B1 (
    .I(MUX_SB_T1_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .O(REG_T1_NORTH_B1_O),
    .CLK(clk),
    .CE(and1_inst4_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T1_SOUTH_B1 (
    .I(MUX_SB_T1_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .O(REG_T1_SOUTH_B1_O),
    .CLK(clk),
    .CE(and1_inst5_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T1_WEST_B1 (
    .I(MUX_SB_T1_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .O(REG_T1_WEST_B1_O),
    .CLK(clk),
    .CE(and1_inst7_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T2_EAST_B1 (
    .I(MUX_SB_T2_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .O(REG_T2_EAST_B1_O),
    .CLK(clk),
    .CE(and1_inst10_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T2_NORTH_B1 (
    .I(MUX_SB_T2_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .O(REG_T2_NORTH_B1_O),
    .CLK(clk),
    .CE(and1_inst8_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T2_SOUTH_B1 (
    .I(MUX_SB_T2_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .O(REG_T2_SOUTH_B1_O),
    .CLK(clk),
    .CE(and1_inst9_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T2_WEST_B1 (
    .I(MUX_SB_T2_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .O(REG_T2_WEST_B1_O),
    .CLK(clk),
    .CE(and1_inst11_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T3_EAST_B1 (
    .I(MUX_SB_T3_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .O(REG_T3_EAST_B1_O),
    .CLK(clk),
    .CE(and1_inst14_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T3_NORTH_B1 (
    .I(MUX_SB_T3_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .O(REG_T3_NORTH_B1_O),
    .CLK(clk),
    .CE(and1_inst12_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T3_SOUTH_B1 (
    .I(MUX_SB_T3_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .O(REG_T3_SOUTH_B1_O),
    .CLK(clk),
    .CE(and1_inst13_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T3_WEST_B1 (
    .I(MUX_SB_T3_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .O(REG_T3_WEST_B1_O),
    .CLK(clk),
    .CE(and1_inst15_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T4_EAST_B1 (
    .I(MUX_SB_T4_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .O(REG_T4_EAST_B1_O),
    .CLK(clk),
    .CE(and1_inst18_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T4_NORTH_B1 (
    .I(MUX_SB_T4_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .O(REG_T4_NORTH_B1_O),
    .CLK(clk),
    .CE(and1_inst16_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T4_SOUTH_B1 (
    .I(MUX_SB_T4_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .O(REG_T4_SOUTH_B1_O),
    .CLK(clk),
    .CE(and1_inst17_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T4_WEST_B1 (
    .I(MUX_SB_T4_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .O(REG_T4_WEST_B1_O),
    .CLK(clk),
    .CE(and1_inst19_out[0])
);
coreir_mux #(
    .width(1)
) RMUX_T0_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T0_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .in1(REG_T0_EAST_B1_O),
    .sel(RMUX_T0_EAST_B1_sel_inst0_O[0]),
    .out(RMUX_T0_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T0_EAST_B1_sel RMUX_T0_EAST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_EAST_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T0_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T0_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .in1(REG_T0_NORTH_B1_O),
    .sel(RMUX_T0_NORTH_B1_sel_inst0_O[0]),
    .out(RMUX_T0_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T0_NORTH_B1_sel RMUX_T0_NORTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_NORTH_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T0_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T0_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .in1(REG_T0_SOUTH_B1_O),
    .sel(RMUX_T0_SOUTH_B1_sel_inst0_O[0]),
    .out(RMUX_T0_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T0_SOUTH_B1_sel RMUX_T0_SOUTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_SOUTH_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T0_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T0_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .in1(REG_T0_WEST_B1_O),
    .sel(RMUX_T0_WEST_B1_sel_inst0_O[0]),
    .out(RMUX_T0_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T0_WEST_B1_sel RMUX_T0_WEST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_WEST_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T1_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T1_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .in1(REG_T1_EAST_B1_O),
    .sel(RMUX_T1_EAST_B1_sel_inst0_O[0]),
    .out(RMUX_T1_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T1_EAST_B1_sel RMUX_T1_EAST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_EAST_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T1_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T1_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .in1(REG_T1_NORTH_B1_O),
    .sel(RMUX_T1_NORTH_B1_sel_inst0_O[0]),
    .out(RMUX_T1_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T1_NORTH_B1_sel RMUX_T1_NORTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_NORTH_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T1_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T1_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .in1(REG_T1_SOUTH_B1_O),
    .sel(RMUX_T1_SOUTH_B1_sel_inst0_O[0]),
    .out(RMUX_T1_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T1_SOUTH_B1_sel RMUX_T1_SOUTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_SOUTH_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T1_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T1_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .in1(REG_T1_WEST_B1_O),
    .sel(RMUX_T1_WEST_B1_sel_inst0_O[0]),
    .out(RMUX_T1_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T1_WEST_B1_sel RMUX_T1_WEST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_WEST_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T2_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T2_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .in1(REG_T2_EAST_B1_O),
    .sel(RMUX_T2_EAST_B1_sel_inst0_O[0]),
    .out(RMUX_T2_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T2_EAST_B1_sel RMUX_T2_EAST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_EAST_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T2_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T2_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .in1(REG_T2_NORTH_B1_O),
    .sel(RMUX_T2_NORTH_B1_sel_inst0_O[0]),
    .out(RMUX_T2_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T2_NORTH_B1_sel RMUX_T2_NORTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_NORTH_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T2_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T2_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .in1(REG_T2_SOUTH_B1_O),
    .sel(RMUX_T2_SOUTH_B1_sel_inst0_O[0]),
    .out(RMUX_T2_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T2_SOUTH_B1_sel RMUX_T2_SOUTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_SOUTH_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T2_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T2_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .in1(REG_T2_WEST_B1_O),
    .sel(RMUX_T2_WEST_B1_sel_inst0_O[0]),
    .out(RMUX_T2_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T2_WEST_B1_sel RMUX_T2_WEST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_WEST_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T3_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T3_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .in1(REG_T3_EAST_B1_O),
    .sel(RMUX_T3_EAST_B1_sel_inst0_O[0]),
    .out(RMUX_T3_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T3_EAST_B1_sel RMUX_T3_EAST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_EAST_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T3_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T3_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .in1(REG_T3_NORTH_B1_O),
    .sel(RMUX_T3_NORTH_B1_sel_inst0_O[0]),
    .out(RMUX_T3_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T3_NORTH_B1_sel RMUX_T3_NORTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_NORTH_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T3_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T3_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .in1(REG_T3_SOUTH_B1_O),
    .sel(RMUX_T3_SOUTH_B1_sel_inst0_O[0]),
    .out(RMUX_T3_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T3_SOUTH_B1_sel RMUX_T3_SOUTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_SOUTH_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T3_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T3_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .in1(REG_T3_WEST_B1_O),
    .sel(RMUX_T3_WEST_B1_sel_inst0_O[0]),
    .out(RMUX_T3_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T3_WEST_B1_sel RMUX_T3_WEST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_WEST_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T4_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T4_EAST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .in1(REG_T4_EAST_B1_O),
    .sel(RMUX_T4_EAST_B1_sel_inst0_O[0]),
    .out(RMUX_T4_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T4_EAST_B1_sel RMUX_T4_EAST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_EAST_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T4_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T4_NORTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .in1(REG_T4_NORTH_B1_O),
    .sel(RMUX_T4_NORTH_B1_sel_inst0_O[0]),
    .out(RMUX_T4_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T4_NORTH_B1_sel RMUX_T4_NORTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_NORTH_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T4_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T4_SOUTH_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .in1(REG_T4_SOUTH_B1_O),
    .sel(RMUX_T4_SOUTH_B1_sel_inst0_O[0]),
    .out(RMUX_T4_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T4_SOUTH_B1_sel RMUX_T4_SOUTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_SOUTH_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T4_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T4_WEST_SB_OUT_B1$Mux9x1_inst0$coreir_commonlib_mux9x1_inst0_out),
    .in1(REG_T4_WEST_B1_O),
    .sel(RMUX_T4_WEST_B1_sel_inst0_O[0]),
    .out(RMUX_T4_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T4_WEST_B1_sel RMUX_T4_WEST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_WEST_B1_sel_inst0_O)
);
SB_T0_EAST_SB_OUT_B1_sel_unq1 SB_T0_EAST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_EAST_SB_OUT_B1_sel_inst0_O)
);
SB_T0_NORTH_SB_OUT_B1_sel_unq1 SB_T0_NORTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_NORTH_SB_OUT_B1_sel_inst0_O)
);
SB_T0_SOUTH_SB_OUT_B1_sel_unq1 SB_T0_SOUTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_SOUTH_SB_OUT_B1_sel_inst0_O)
);
SB_T0_WEST_SB_OUT_B1_sel_unq1 SB_T0_WEST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T0_WEST_SB_OUT_B1_sel_inst0_O)
);
SB_T1_EAST_SB_OUT_B1_sel_unq1 SB_T1_EAST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_EAST_SB_OUT_B1_sel_inst0_O)
);
SB_T1_NORTH_SB_OUT_B1_sel_unq1 SB_T1_NORTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_NORTH_SB_OUT_B1_sel_inst0_O)
);
SB_T1_SOUTH_SB_OUT_B1_sel_unq1 SB_T1_SOUTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_SOUTH_SB_OUT_B1_sel_inst0_O)
);
SB_T1_WEST_SB_OUT_B1_sel_unq1 SB_T1_WEST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_WEST_SB_OUT_B1_sel_inst0_O)
);
SB_T2_EAST_SB_OUT_B1_sel_unq1 SB_T2_EAST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_EAST_SB_OUT_B1_sel_inst0_O)
);
SB_T2_NORTH_SB_OUT_B1_sel_unq1 SB_T2_NORTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_NORTH_SB_OUT_B1_sel_inst0_O)
);
SB_T2_SOUTH_SB_OUT_B1_sel_unq1 SB_T2_SOUTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_SOUTH_SB_OUT_B1_sel_inst0_O)
);
SB_T2_WEST_SB_OUT_B1_sel_unq1 SB_T2_WEST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T2_WEST_SB_OUT_B1_sel_inst0_O)
);
SB_T3_EAST_SB_OUT_B1_sel_unq1 SB_T3_EAST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T3_EAST_SB_OUT_B1_sel_inst0_O)
);
SB_T3_NORTH_SB_OUT_B1_sel_unq1 SB_T3_NORTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T3_NORTH_SB_OUT_B1_sel_inst0_O)
);
SB_T3_SOUTH_SB_OUT_B1_sel_unq1 SB_T3_SOUTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T3_SOUTH_SB_OUT_B1_sel_inst0_O)
);
SB_T3_WEST_SB_OUT_B1_sel_unq1 SB_T3_WEST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T3_WEST_SB_OUT_B1_sel_inst0_O)
);
SB_T4_EAST_SB_OUT_B1_sel_unq1 SB_T4_EAST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T4_EAST_SB_OUT_B1_sel_inst0_O)
);
SB_T4_NORTH_SB_OUT_B1_sel_unq1 SB_T4_NORTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T4_NORTH_SB_OUT_B1_sel_inst0_O)
);
SB_T4_SOUTH_SB_OUT_B1_sel_unq1 SB_T4_SOUTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T4_SOUTH_SB_OUT_B1_sel_inst0_O)
);
SB_T4_WEST_SB_OUT_B1_sel_unq1 SB_T4_WEST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_3_O),
    .O(SB_T4_WEST_SB_OUT_B1_sel_inst0_O)
);
MuxWrapper_1_1 WIRE_SB_T0_EAST_SB_IN_B1 (
    .I(SB_T0_EAST_SB_IN_B1),
    .O(WIRE_SB_T0_EAST_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T0_NORTH_SB_IN_B1 (
    .I(SB_T0_NORTH_SB_IN_B1),
    .O(WIRE_SB_T0_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T0_SOUTH_SB_IN_B1 (
    .I(SB_T0_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T0_WEST_SB_IN_B1 (
    .I(SB_T0_WEST_SB_IN_B1),
    .O(WIRE_SB_T0_WEST_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T1_EAST_SB_IN_B1 (
    .I(SB_T1_EAST_SB_IN_B1),
    .O(WIRE_SB_T1_EAST_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T1_NORTH_SB_IN_B1 (
    .I(SB_T1_NORTH_SB_IN_B1),
    .O(WIRE_SB_T1_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T1_SOUTH_SB_IN_B1 (
    .I(SB_T1_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T1_WEST_SB_IN_B1 (
    .I(SB_T1_WEST_SB_IN_B1),
    .O(WIRE_SB_T1_WEST_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T2_EAST_SB_IN_B1 (
    .I(SB_T2_EAST_SB_IN_B1),
    .O(WIRE_SB_T2_EAST_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T2_NORTH_SB_IN_B1 (
    .I(SB_T2_NORTH_SB_IN_B1),
    .O(WIRE_SB_T2_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T2_SOUTH_SB_IN_B1 (
    .I(SB_T2_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T2_WEST_SB_IN_B1 (
    .I(SB_T2_WEST_SB_IN_B1),
    .O(WIRE_SB_T2_WEST_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T3_EAST_SB_IN_B1 (
    .I(SB_T3_EAST_SB_IN_B1),
    .O(WIRE_SB_T3_EAST_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T3_NORTH_SB_IN_B1 (
    .I(SB_T3_NORTH_SB_IN_B1),
    .O(WIRE_SB_T3_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T3_SOUTH_SB_IN_B1 (
    .I(SB_T3_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T3_WEST_SB_IN_B1 (
    .I(SB_T3_WEST_SB_IN_B1),
    .O(WIRE_SB_T3_WEST_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T4_EAST_SB_IN_B1 (
    .I(SB_T4_EAST_SB_IN_B1),
    .O(WIRE_SB_T4_EAST_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T4_NORTH_SB_IN_B1 (
    .I(SB_T4_NORTH_SB_IN_B1),
    .O(WIRE_SB_T4_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T4_SOUTH_SB_IN_B1 (
    .I(SB_T4_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T4_WEST_SB_IN_B1 (
    .I(SB_T4_WEST_SB_IN_B1),
    .O(WIRE_SB_T4_WEST_SB_IN_B1_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_4_32_inst0$bit_const_0_None (
    .out(ZextWrapper_4_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit4 ZextWrapper_4_32_inst0$self_I (
    .in(config_reg_3_O),
    .out(ZextWrapper_4_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_4_32_inst0$self_O_out;
assign ZextWrapper_4_32_inst0$self_O_out = {ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$bit_const_0_None_out,ZextWrapper_4_32_inst0$self_I_out[3:0]};
mantle_wire__typeBitIn32 ZextWrapper_4_32_inst0$self_O (
    .in(ZextWrapper_4_32_inst0$self_O_in),
    .out(ZextWrapper_4_32_inst0$self_O_out)
);
coreir_and #(
    .width(1)
) and1_inst0 (
    .in0(coreir_eq_1_inst0_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst0_out)
);
coreir_and #(
    .width(1)
) and1_inst1 (
    .in0(coreir_eq_1_inst1_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst1_out)
);
coreir_and #(
    .width(1)
) and1_inst10 (
    .in0(coreir_eq_1_inst10_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst10_out)
);
coreir_and #(
    .width(1)
) and1_inst11 (
    .in0(coreir_eq_1_inst11_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst11_out)
);
coreir_and #(
    .width(1)
) and1_inst12 (
    .in0(coreir_eq_1_inst12_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst12_out)
);
coreir_and #(
    .width(1)
) and1_inst13 (
    .in0(coreir_eq_1_inst13_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst13_out)
);
coreir_and #(
    .width(1)
) and1_inst14 (
    .in0(coreir_eq_1_inst14_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst14_out)
);
coreir_and #(
    .width(1)
) and1_inst15 (
    .in0(coreir_eq_1_inst15_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst15_out)
);
coreir_and #(
    .width(1)
) and1_inst16 (
    .in0(coreir_eq_1_inst16_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst16_out)
);
coreir_and #(
    .width(1)
) and1_inst17 (
    .in0(coreir_eq_1_inst17_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst17_out)
);
coreir_and #(
    .width(1)
) and1_inst18 (
    .in0(coreir_eq_1_inst18_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst18_out)
);
coreir_and #(
    .width(1)
) and1_inst19 (
    .in0(coreir_eq_1_inst19_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst19_out)
);
coreir_and #(
    .width(1)
) and1_inst2 (
    .in0(coreir_eq_1_inst2_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst2_out)
);
coreir_and #(
    .width(1)
) and1_inst3 (
    .in0(coreir_eq_1_inst3_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst3_out)
);
coreir_and #(
    .width(1)
) and1_inst4 (
    .in0(coreir_eq_1_inst4_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst4_out)
);
coreir_and #(
    .width(1)
) and1_inst5 (
    .in0(coreir_eq_1_inst5_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst5_out)
);
coreir_and #(
    .width(1)
) and1_inst6 (
    .in0(coreir_eq_1_inst6_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst6_out)
);
coreir_and #(
    .width(1)
) and1_inst7 (
    .in0(coreir_eq_1_inst7_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst7_out)
);
coreir_and #(
    .width(1)
) and1_inst8 (
    .in0(coreir_eq_1_inst8_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst8_out)
);
coreir_and #(
    .width(1)
) and1_inst9 (
    .in0(coreir_eq_1_inst9_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst9_out)
);
ConfigRegister_32_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_1 config_reg_1 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_1_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_2 config_reg_2 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_2_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_4_8_32_3 config_reg_3 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_3_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
coreir_const #(
    .value(1'h1),
    .width(1)
) const_1_1 (
    .out(const_1_1_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst0 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_NORTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst0_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst1 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_SOUTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst1_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst10 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_EAST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst10_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst11 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_WEST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst11_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst12 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_NORTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst12_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst13 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_SOUTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst13_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst14 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_EAST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst14_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst15 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_WEST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst15_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst16 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_NORTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst16_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst17 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_SOUTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst17_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst18 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_EAST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst18_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst19 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_WEST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst19_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst2 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_EAST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst2_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst3 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_WEST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst3_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst4 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_NORTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst4_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst5 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_SOUTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst5_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst6 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_EAST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst6_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst7 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_WEST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst7_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst8 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_NORTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst8_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst9 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_SOUTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst9_out)
);
mantle_wire__typeBit8 self_config_config_addr (
    .in(config_config_addr),
    .out(self_config_config_addr_out)
);
assign SB_T0_EAST_SB_OUT_B1 = RMUX_T0_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T0_NORTH_SB_OUT_B1 = RMUX_T0_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T0_SOUTH_SB_OUT_B1 = RMUX_T0_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T0_WEST_SB_OUT_B1 = RMUX_T0_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T1_EAST_SB_OUT_B1 = RMUX_T1_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T1_NORTH_SB_OUT_B1 = RMUX_T1_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T1_SOUTH_SB_OUT_B1 = RMUX_T1_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T1_WEST_SB_OUT_B1 = RMUX_T1_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T2_EAST_SB_OUT_B1 = RMUX_T2_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T2_NORTH_SB_OUT_B1 = RMUX_T2_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T2_SOUTH_SB_OUT_B1 = RMUX_T2_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T2_WEST_SB_OUT_B1 = RMUX_T2_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T3_EAST_SB_OUT_B1 = RMUX_T3_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T3_NORTH_SB_OUT_B1 = RMUX_T3_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T3_SOUTH_SB_OUT_B1 = RMUX_T3_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T3_WEST_SB_OUT_B1 = RMUX_T3_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T4_EAST_SB_OUT_B1 = RMUX_T4_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T4_NORTH_SB_OUT_B1 = RMUX_T4_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T4_SOUTH_SB_OUT_B1 = RMUX_T4_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T4_WEST_SB_OUT_B1 = RMUX_T4_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign read_config_data = MuxWrapper_4_32_inst0$Mux4x32_inst0$coreir_commonlib_mux4x32_inst0_out;
endmodule

module ConfigRegister_31_8_32_50 (
    input clk,
    input reset,
    output [30:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [30:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_31_inst0_O;
wire [7:0] const_50_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_31 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_31_inst0 (
    .I(config_data[30:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_31_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h32),
    .width(8)
) const_50_8 (
    .out(const_50_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_50_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_31_inst0_O;
endmodule

module ConfigRegister_30_8_32_1 (
    input clk,
    input reset,
    output [29:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [29:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_30_inst0_O;
wire [7:0] const_1_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_30 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_30_inst0 (
    .I(config_data[29:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_30_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h01),
    .width(8)
) const_1_8 (
    .out(const_1_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_1_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_30_inst0_O;
endmodule

module ConfigRegister_29_8_32_83 (
    input clk,
    input reset,
    output [28:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [28:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_29_inst0_O;
wire [7:0] const_83_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_29 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_29_inst0 (
    .I(config_data[28:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_29_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h53),
    .width(8)
) const_83_8 (
    .out(const_83_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_83_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_29_inst0_O;
endmodule

module ConfigRegister_28_8_32_1 (
    input clk,
    input reset,
    output [27:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [27:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_28_inst0_O;
wire [7:0] const_1_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_28 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_28_inst0 (
    .I(config_data[27:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_28_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h01),
    .width(8)
) const_1_8 (
    .out(const_1_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_1_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_28_inst0_O;
endmodule

module SB_ID0_5TRACKS_B1_PE (
    input [0:0] SB_T0_EAST_SB_IN_B1,
    output [0:0] SB_T0_EAST_SB_OUT_B1,
    input [0:0] SB_T0_NORTH_SB_IN_B1,
    output [0:0] SB_T0_NORTH_SB_OUT_B1,
    input [0:0] SB_T0_SOUTH_SB_IN_B1,
    output [0:0] SB_T0_SOUTH_SB_OUT_B1,
    input [0:0] SB_T0_WEST_SB_IN_B1,
    output [0:0] SB_T0_WEST_SB_OUT_B1,
    input [0:0] SB_T1_EAST_SB_IN_B1,
    output [0:0] SB_T1_EAST_SB_OUT_B1,
    input [0:0] SB_T1_NORTH_SB_IN_B1,
    output [0:0] SB_T1_NORTH_SB_OUT_B1,
    input [0:0] SB_T1_SOUTH_SB_IN_B1,
    output [0:0] SB_T1_SOUTH_SB_OUT_B1,
    input [0:0] SB_T1_WEST_SB_IN_B1,
    output [0:0] SB_T1_WEST_SB_OUT_B1,
    input [0:0] SB_T2_EAST_SB_IN_B1,
    output [0:0] SB_T2_EAST_SB_OUT_B1,
    input [0:0] SB_T2_NORTH_SB_IN_B1,
    output [0:0] SB_T2_NORTH_SB_OUT_B1,
    input [0:0] SB_T2_SOUTH_SB_IN_B1,
    output [0:0] SB_T2_SOUTH_SB_OUT_B1,
    input [0:0] SB_T2_WEST_SB_IN_B1,
    output [0:0] SB_T2_WEST_SB_OUT_B1,
    input [0:0] SB_T3_EAST_SB_IN_B1,
    output [0:0] SB_T3_EAST_SB_OUT_B1,
    input [0:0] SB_T3_NORTH_SB_IN_B1,
    output [0:0] SB_T3_NORTH_SB_OUT_B1,
    input [0:0] SB_T3_SOUTH_SB_IN_B1,
    output [0:0] SB_T3_SOUTH_SB_OUT_B1,
    input [0:0] SB_T3_WEST_SB_IN_B1,
    output [0:0] SB_T3_WEST_SB_OUT_B1,
    input [0:0] SB_T4_EAST_SB_IN_B1,
    output [0:0] SB_T4_EAST_SB_OUT_B1,
    input [0:0] SB_T4_NORTH_SB_IN_B1,
    output [0:0] SB_T4_NORTH_SB_OUT_B1,
    input [0:0] SB_T4_SOUTH_SB_IN_B1,
    output [0:0] SB_T4_SOUTH_SB_OUT_B1,
    input [0:0] SB_T4_WEST_SB_IN_B1,
    output [0:0] SB_T4_WEST_SB_OUT_B1,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    input [0:0] pe_outputs_1,
    output [31:0] read_config_data,
    input reset,
    input [0:0] stall
);
wire [0:0] Invert1_inst0_out;
wire [0:0] MUX_SB_T0_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out;
wire [0:0] MUX_SB_T0_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out;
wire [0:0] MUX_SB_T0_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out;
wire [0:0] MUX_SB_T0_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out;
wire [0:0] MUX_SB_T1_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out;
wire [0:0] MUX_SB_T1_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out;
wire [0:0] MUX_SB_T1_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out;
wire [0:0] MUX_SB_T1_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out;
wire [0:0] MUX_SB_T2_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out;
wire [0:0] MUX_SB_T2_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out;
wire [0:0] MUX_SB_T2_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out;
wire [0:0] MUX_SB_T2_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out;
wire [0:0] MUX_SB_T3_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out;
wire [0:0] MUX_SB_T3_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out;
wire [0:0] MUX_SB_T3_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out;
wire [0:0] MUX_SB_T3_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out;
wire [0:0] MUX_SB_T4_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out;
wire [0:0] MUX_SB_T4_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out;
wire [0:0] MUX_SB_T4_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out;
wire [0:0] MUX_SB_T4_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out;
wire [31:0] MuxWrapper_2_32_inst0$Mux2x32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
wire [0:0] REG_T0_EAST_B1_O;
wire [0:0] REG_T0_NORTH_B1_O;
wire [0:0] REG_T0_SOUTH_B1_O;
wire [0:0] REG_T0_WEST_B1_O;
wire [0:0] REG_T1_EAST_B1_O;
wire [0:0] REG_T1_NORTH_B1_O;
wire [0:0] REG_T1_SOUTH_B1_O;
wire [0:0] REG_T1_WEST_B1_O;
wire [0:0] REG_T2_EAST_B1_O;
wire [0:0] REG_T2_NORTH_B1_O;
wire [0:0] REG_T2_SOUTH_B1_O;
wire [0:0] REG_T2_WEST_B1_O;
wire [0:0] REG_T3_EAST_B1_O;
wire [0:0] REG_T3_NORTH_B1_O;
wire [0:0] REG_T3_SOUTH_B1_O;
wire [0:0] REG_T3_WEST_B1_O;
wire [0:0] REG_T4_EAST_B1_O;
wire [0:0] REG_T4_NORTH_B1_O;
wire [0:0] REG_T4_SOUTH_B1_O;
wire [0:0] REG_T4_WEST_B1_O;
wire [0:0] RMUX_T0_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T0_EAST_B1_sel_inst0_O;
wire [0:0] RMUX_T0_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T0_NORTH_B1_sel_inst0_O;
wire [0:0] RMUX_T0_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T0_SOUTH_B1_sel_inst0_O;
wire [0:0] RMUX_T0_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T0_WEST_B1_sel_inst0_O;
wire [0:0] RMUX_T1_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T1_EAST_B1_sel_inst0_O;
wire [0:0] RMUX_T1_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T1_NORTH_B1_sel_inst0_O;
wire [0:0] RMUX_T1_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T1_SOUTH_B1_sel_inst0_O;
wire [0:0] RMUX_T1_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T1_WEST_B1_sel_inst0_O;
wire [0:0] RMUX_T2_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T2_EAST_B1_sel_inst0_O;
wire [0:0] RMUX_T2_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T2_NORTH_B1_sel_inst0_O;
wire [0:0] RMUX_T2_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T2_SOUTH_B1_sel_inst0_O;
wire [0:0] RMUX_T2_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T2_WEST_B1_sel_inst0_O;
wire [0:0] RMUX_T3_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T3_EAST_B1_sel_inst0_O;
wire [0:0] RMUX_T3_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T3_NORTH_B1_sel_inst0_O;
wire [0:0] RMUX_T3_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T3_SOUTH_B1_sel_inst0_O;
wire [0:0] RMUX_T3_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T3_WEST_B1_sel_inst0_O;
wire [0:0] RMUX_T4_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T4_EAST_B1_sel_inst0_O;
wire [0:0] RMUX_T4_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T4_NORTH_B1_sel_inst0_O;
wire [0:0] RMUX_T4_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T4_SOUTH_B1_sel_inst0_O;
wire [0:0] RMUX_T4_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] RMUX_T4_WEST_B1_sel_inst0_O;
wire [1:0] SB_T0_EAST_SB_OUT_B1_sel_inst0_O;
wire [1:0] SB_T0_NORTH_SB_OUT_B1_sel_inst0_O;
wire [1:0] SB_T0_SOUTH_SB_OUT_B1_sel_inst0_O;
wire [1:0] SB_T0_WEST_SB_OUT_B1_sel_inst0_O;
wire [1:0] SB_T1_EAST_SB_OUT_B1_sel_inst0_O;
wire [1:0] SB_T1_NORTH_SB_OUT_B1_sel_inst0_O;
wire [1:0] SB_T1_SOUTH_SB_OUT_B1_sel_inst0_O;
wire [1:0] SB_T1_WEST_SB_OUT_B1_sel_inst0_O;
wire [1:0] SB_T2_EAST_SB_OUT_B1_sel_inst0_O;
wire [1:0] SB_T2_NORTH_SB_OUT_B1_sel_inst0_O;
wire [1:0] SB_T2_SOUTH_SB_OUT_B1_sel_inst0_O;
wire [1:0] SB_T2_WEST_SB_OUT_B1_sel_inst0_O;
wire [1:0] SB_T3_EAST_SB_OUT_B1_sel_inst0_O;
wire [1:0] SB_T3_NORTH_SB_OUT_B1_sel_inst0_O;
wire [1:0] SB_T3_SOUTH_SB_OUT_B1_sel_inst0_O;
wire [1:0] SB_T3_WEST_SB_OUT_B1_sel_inst0_O;
wire [1:0] SB_T4_EAST_SB_OUT_B1_sel_inst0_O;
wire [1:0] SB_T4_NORTH_SB_OUT_B1_sel_inst0_O;
wire [1:0] SB_T4_SOUTH_SB_OUT_B1_sel_inst0_O;
wire [1:0] SB_T4_WEST_SB_OUT_B1_sel_inst0_O;
wire [0:0] WIRE_SB_T0_EAST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T0_NORTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T0_SOUTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T0_WEST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T1_EAST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T1_NORTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T1_SOUTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T1_WEST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T2_EAST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T2_NORTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T2_SOUTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T2_WEST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T3_EAST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T3_NORTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T3_SOUTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T3_WEST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T4_EAST_SB_IN_B1_O;
wire [0:0] WIRE_SB_T4_NORTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T4_SOUTH_SB_IN_B1_O;
wire [0:0] WIRE_SB_T4_WEST_SB_IN_B1_O;
wire ZextWrapper_28_32_inst0$bit_const_0_None_out;
wire [27:0] ZextWrapper_28_32_inst0$self_I_out;
wire [31:0] ZextWrapper_28_32_inst0$self_O_in;
wire [0:0] and1_inst0_out;
wire [0:0] and1_inst1_out;
wire [0:0] and1_inst10_out;
wire [0:0] and1_inst11_out;
wire [0:0] and1_inst12_out;
wire [0:0] and1_inst13_out;
wire [0:0] and1_inst14_out;
wire [0:0] and1_inst15_out;
wire [0:0] and1_inst16_out;
wire [0:0] and1_inst17_out;
wire [0:0] and1_inst18_out;
wire [0:0] and1_inst19_out;
wire [0:0] and1_inst2_out;
wire [0:0] and1_inst3_out;
wire [0:0] and1_inst4_out;
wire [0:0] and1_inst5_out;
wire [0:0] and1_inst6_out;
wire [0:0] and1_inst7_out;
wire [0:0] and1_inst8_out;
wire [0:0] and1_inst9_out;
wire [31:0] config_reg_0_O;
wire [27:0] config_reg_1_O;
wire [0:0] const_1_1_out;
wire coreir_eq_1_inst0_out;
wire coreir_eq_1_inst1_out;
wire coreir_eq_1_inst10_out;
wire coreir_eq_1_inst11_out;
wire coreir_eq_1_inst12_out;
wire coreir_eq_1_inst13_out;
wire coreir_eq_1_inst14_out;
wire coreir_eq_1_inst15_out;
wire coreir_eq_1_inst16_out;
wire coreir_eq_1_inst17_out;
wire coreir_eq_1_inst18_out;
wire coreir_eq_1_inst19_out;
wire coreir_eq_1_inst2_out;
wire coreir_eq_1_inst3_out;
wire coreir_eq_1_inst4_out;
wire coreir_eq_1_inst5_out;
wire coreir_eq_1_inst6_out;
wire coreir_eq_1_inst7_out;
wire coreir_eq_1_inst8_out;
wire coreir_eq_1_inst9_out;
coreir_not #(
    .width(1)
) Invert1_inst0 (
    .in(stall),
    .out(Invert1_inst0_out)
);
commonlib_muxn__N4__width1 MUX_SB_T0_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0 (
    .in_data_0(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .in_data_3(pe_outputs_1),
    .in_sel(SB_T0_EAST_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T0_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out)
);
commonlib_muxn__N4__width1 MUX_SB_T0_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0 (
    .in_data_0(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .in_data_3(pe_outputs_1),
    .in_sel(SB_T0_NORTH_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T0_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out)
);
commonlib_muxn__N4__width1 MUX_SB_T0_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0 (
    .in_data_0(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .in_data_3(pe_outputs_1),
    .in_sel(SB_T0_SOUTH_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T0_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out)
);
commonlib_muxn__N4__width1 MUX_SB_T0_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0 (
    .in_data_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .in_data_3(pe_outputs_1),
    .in_sel(SB_T0_WEST_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T0_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out)
);
commonlib_muxn__N4__width1 MUX_SB_T1_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0 (
    .in_data_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .in_data_3(pe_outputs_1),
    .in_sel(SB_T1_EAST_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T1_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out)
);
commonlib_muxn__N4__width1 MUX_SB_T1_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0 (
    .in_data_0(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .in_data_3(pe_outputs_1),
    .in_sel(SB_T1_NORTH_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T1_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out)
);
commonlib_muxn__N4__width1 MUX_SB_T1_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0 (
    .in_data_0(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .in_data_3(pe_outputs_1),
    .in_sel(SB_T1_SOUTH_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T1_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out)
);
commonlib_muxn__N4__width1 MUX_SB_T1_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0 (
    .in_data_0(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .in_data_3(pe_outputs_1),
    .in_sel(SB_T1_WEST_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T1_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out)
);
commonlib_muxn__N4__width1 MUX_SB_T2_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0 (
    .in_data_0(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .in_data_3(pe_outputs_1),
    .in_sel(SB_T2_EAST_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T2_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out)
);
commonlib_muxn__N4__width1 MUX_SB_T2_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0 (
    .in_data_0(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .in_data_3(pe_outputs_1),
    .in_sel(SB_T2_NORTH_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T2_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out)
);
commonlib_muxn__N4__width1 MUX_SB_T2_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0 (
    .in_data_0(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .in_data_3(pe_outputs_1),
    .in_sel(SB_T2_SOUTH_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T2_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out)
);
commonlib_muxn__N4__width1 MUX_SB_T2_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0 (
    .in_data_0(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .in_data_3(pe_outputs_1),
    .in_sel(SB_T2_WEST_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T2_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out)
);
commonlib_muxn__N4__width1 MUX_SB_T3_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0 (
    .in_data_0(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .in_data_3(pe_outputs_1),
    .in_sel(SB_T3_EAST_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T3_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out)
);
commonlib_muxn__N4__width1 MUX_SB_T3_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0 (
    .in_data_0(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .in_data_3(pe_outputs_1),
    .in_sel(SB_T3_NORTH_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T3_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out)
);
commonlib_muxn__N4__width1 MUX_SB_T3_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0 (
    .in_data_0(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .in_data_3(pe_outputs_1),
    .in_sel(SB_T3_SOUTH_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T3_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out)
);
commonlib_muxn__N4__width1 MUX_SB_T3_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0 (
    .in_data_0(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .in_data_3(pe_outputs_1),
    .in_sel(SB_T3_WEST_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T3_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out)
);
commonlib_muxn__N4__width1 MUX_SB_T4_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0 (
    .in_data_0(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .in_data_3(pe_outputs_1),
    .in_sel(SB_T4_EAST_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T4_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out)
);
commonlib_muxn__N4__width1 MUX_SB_T4_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0 (
    .in_data_0(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .in_data_3(pe_outputs_1),
    .in_sel(SB_T4_NORTH_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T4_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out)
);
commonlib_muxn__N4__width1 MUX_SB_T4_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0 (
    .in_data_0(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .in_data_3(pe_outputs_1),
    .in_sel(SB_T4_SOUTH_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T4_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out)
);
commonlib_muxn__N4__width1 MUX_SB_T4_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0 (
    .in_data_0(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .in_data_1(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .in_data_2(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .in_data_3(pe_outputs_1),
    .in_sel(SB_T4_WEST_SB_OUT_B1_sel_inst0_O),
    .out(MUX_SB_T4_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out)
);
coreir_mux #(
    .width(32)
) MuxWrapper_2_32_inst0$Mux2x32_inst0$coreir_commonlib_mux2x32_inst0$_join (
    .in0(config_reg_0_O),
    .in1(ZextWrapper_28_32_inst0$self_O_in),
    .sel(config_config_addr[0]),
    .out(MuxWrapper_2_32_inst0$Mux2x32_inst0$coreir_commonlib_mux2x32_inst0$_join_out)
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T0_EAST_B1 (
    .I(MUX_SB_T0_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .O(REG_T0_EAST_B1_O),
    .CLK(clk),
    .CE(and1_inst2_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T0_NORTH_B1 (
    .I(MUX_SB_T0_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .O(REG_T0_NORTH_B1_O),
    .CLK(clk),
    .CE(and1_inst0_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T0_SOUTH_B1 (
    .I(MUX_SB_T0_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .O(REG_T0_SOUTH_B1_O),
    .CLK(clk),
    .CE(and1_inst1_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T0_WEST_B1 (
    .I(MUX_SB_T0_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .O(REG_T0_WEST_B1_O),
    .CLK(clk),
    .CE(and1_inst3_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T1_EAST_B1 (
    .I(MUX_SB_T1_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .O(REG_T1_EAST_B1_O),
    .CLK(clk),
    .CE(and1_inst6_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T1_NORTH_B1 (
    .I(MUX_SB_T1_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .O(REG_T1_NORTH_B1_O),
    .CLK(clk),
    .CE(and1_inst4_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T1_SOUTH_B1 (
    .I(MUX_SB_T1_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .O(REG_T1_SOUTH_B1_O),
    .CLK(clk),
    .CE(and1_inst5_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T1_WEST_B1 (
    .I(MUX_SB_T1_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .O(REG_T1_WEST_B1_O),
    .CLK(clk),
    .CE(and1_inst7_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T2_EAST_B1 (
    .I(MUX_SB_T2_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .O(REG_T2_EAST_B1_O),
    .CLK(clk),
    .CE(and1_inst10_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T2_NORTH_B1 (
    .I(MUX_SB_T2_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .O(REG_T2_NORTH_B1_O),
    .CLK(clk),
    .CE(and1_inst8_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T2_SOUTH_B1 (
    .I(MUX_SB_T2_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .O(REG_T2_SOUTH_B1_O),
    .CLK(clk),
    .CE(and1_inst9_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T2_WEST_B1 (
    .I(MUX_SB_T2_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .O(REG_T2_WEST_B1_O),
    .CLK(clk),
    .CE(and1_inst11_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T3_EAST_B1 (
    .I(MUX_SB_T3_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .O(REG_T3_EAST_B1_O),
    .CLK(clk),
    .CE(and1_inst14_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T3_NORTH_B1 (
    .I(MUX_SB_T3_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .O(REG_T3_NORTH_B1_O),
    .CLK(clk),
    .CE(and1_inst12_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T3_SOUTH_B1 (
    .I(MUX_SB_T3_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .O(REG_T3_SOUTH_B1_O),
    .CLK(clk),
    .CE(and1_inst13_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T3_WEST_B1 (
    .I(MUX_SB_T3_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .O(REG_T3_WEST_B1_O),
    .CLK(clk),
    .CE(and1_inst15_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T4_EAST_B1 (
    .I(MUX_SB_T4_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .O(REG_T4_EAST_B1_O),
    .CLK(clk),
    .CE(and1_inst18_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T4_NORTH_B1 (
    .I(MUX_SB_T4_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .O(REG_T4_NORTH_B1_O),
    .CLK(clk),
    .CE(and1_inst16_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T4_SOUTH_B1 (
    .I(MUX_SB_T4_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .O(REG_T4_SOUTH_B1_O),
    .CLK(clk),
    .CE(and1_inst17_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_1 REG_T4_WEST_B1 (
    .I(MUX_SB_T4_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .O(REG_T4_WEST_B1_O),
    .CLK(clk),
    .CE(and1_inst19_out[0])
);
coreir_mux #(
    .width(1)
) RMUX_T0_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T0_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .in1(REG_T0_EAST_B1_O),
    .sel(RMUX_T0_EAST_B1_sel_inst0_O[0]),
    .out(RMUX_T0_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T0_EAST_B1_sel RMUX_T0_EAST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_EAST_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T0_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T0_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .in1(REG_T0_NORTH_B1_O),
    .sel(RMUX_T0_NORTH_B1_sel_inst0_O[0]),
    .out(RMUX_T0_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T0_NORTH_B1_sel RMUX_T0_NORTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_NORTH_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T0_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T0_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .in1(REG_T0_SOUTH_B1_O),
    .sel(RMUX_T0_SOUTH_B1_sel_inst0_O[0]),
    .out(RMUX_T0_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T0_SOUTH_B1_sel RMUX_T0_SOUTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_SOUTH_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T0_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T0_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .in1(REG_T0_WEST_B1_O),
    .sel(RMUX_T0_WEST_B1_sel_inst0_O[0]),
    .out(RMUX_T0_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T0_WEST_B1_sel RMUX_T0_WEST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_WEST_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T1_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T1_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .in1(REG_T1_EAST_B1_O),
    .sel(RMUX_T1_EAST_B1_sel_inst0_O[0]),
    .out(RMUX_T1_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T1_EAST_B1_sel RMUX_T1_EAST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_EAST_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T1_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T1_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .in1(REG_T1_NORTH_B1_O),
    .sel(RMUX_T1_NORTH_B1_sel_inst0_O[0]),
    .out(RMUX_T1_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T1_NORTH_B1_sel RMUX_T1_NORTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_NORTH_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T1_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T1_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .in1(REG_T1_SOUTH_B1_O),
    .sel(RMUX_T1_SOUTH_B1_sel_inst0_O[0]),
    .out(RMUX_T1_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T1_SOUTH_B1_sel RMUX_T1_SOUTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_SOUTH_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T1_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T1_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .in1(REG_T1_WEST_B1_O),
    .sel(RMUX_T1_WEST_B1_sel_inst0_O[0]),
    .out(RMUX_T1_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T1_WEST_B1_sel RMUX_T1_WEST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_WEST_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T2_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T2_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .in1(REG_T2_EAST_B1_O),
    .sel(RMUX_T2_EAST_B1_sel_inst0_O[0]),
    .out(RMUX_T2_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T2_EAST_B1_sel RMUX_T2_EAST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_EAST_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T2_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T2_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .in1(REG_T2_NORTH_B1_O),
    .sel(RMUX_T2_NORTH_B1_sel_inst0_O[0]),
    .out(RMUX_T2_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T2_NORTH_B1_sel RMUX_T2_NORTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_NORTH_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T2_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T2_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .in1(REG_T2_SOUTH_B1_O),
    .sel(RMUX_T2_SOUTH_B1_sel_inst0_O[0]),
    .out(RMUX_T2_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T2_SOUTH_B1_sel RMUX_T2_SOUTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_SOUTH_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T2_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T2_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .in1(REG_T2_WEST_B1_O),
    .sel(RMUX_T2_WEST_B1_sel_inst0_O[0]),
    .out(RMUX_T2_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T2_WEST_B1_sel RMUX_T2_WEST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_WEST_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T3_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T3_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .in1(REG_T3_EAST_B1_O),
    .sel(RMUX_T3_EAST_B1_sel_inst0_O[0]),
    .out(RMUX_T3_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T3_EAST_B1_sel RMUX_T3_EAST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_EAST_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T3_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T3_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .in1(REG_T3_NORTH_B1_O),
    .sel(RMUX_T3_NORTH_B1_sel_inst0_O[0]),
    .out(RMUX_T3_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T3_NORTH_B1_sel RMUX_T3_NORTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_NORTH_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T3_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T3_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .in1(REG_T3_SOUTH_B1_O),
    .sel(RMUX_T3_SOUTH_B1_sel_inst0_O[0]),
    .out(RMUX_T3_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T3_SOUTH_B1_sel RMUX_T3_SOUTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_SOUTH_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T3_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T3_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .in1(REG_T3_WEST_B1_O),
    .sel(RMUX_T3_WEST_B1_sel_inst0_O[0]),
    .out(RMUX_T3_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T3_WEST_B1_sel RMUX_T3_WEST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_WEST_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T4_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T4_EAST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .in1(REG_T4_EAST_B1_O),
    .sel(RMUX_T4_EAST_B1_sel_inst0_O[0]),
    .out(RMUX_T4_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T4_EAST_B1_sel RMUX_T4_EAST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_EAST_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T4_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T4_NORTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .in1(REG_T4_NORTH_B1_O),
    .sel(RMUX_T4_NORTH_B1_sel_inst0_O[0]),
    .out(RMUX_T4_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T4_NORTH_B1_sel RMUX_T4_NORTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_NORTH_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T4_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T4_SOUTH_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .in1(REG_T4_SOUTH_B1_O),
    .sel(RMUX_T4_SOUTH_B1_sel_inst0_O[0]),
    .out(RMUX_T4_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T4_SOUTH_B1_sel RMUX_T4_SOUTH_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_SOUTH_B1_sel_inst0_O)
);
coreir_mux #(
    .width(1)
) RMUX_T4_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(MUX_SB_T4_WEST_SB_OUT_B1$Mux4x1_inst0$coreir_commonlib_mux4x1_inst0_out),
    .in1(REG_T4_WEST_B1_O),
    .sel(RMUX_T4_WEST_B1_sel_inst0_O[0]),
    .out(RMUX_T4_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
RMUX_T4_WEST_B1_sel RMUX_T4_WEST_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_WEST_B1_sel_inst0_O)
);
SB_T0_EAST_SB_OUT_B1_sel SB_T0_EAST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_EAST_SB_OUT_B1_sel_inst0_O)
);
SB_T0_NORTH_SB_OUT_B1_sel SB_T0_NORTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_NORTH_SB_OUT_B1_sel_inst0_O)
);
SB_T0_SOUTH_SB_OUT_B1_sel SB_T0_SOUTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_SOUTH_SB_OUT_B1_sel_inst0_O)
);
SB_T0_WEST_SB_OUT_B1_sel SB_T0_WEST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_WEST_SB_OUT_B1_sel_inst0_O)
);
SB_T1_EAST_SB_OUT_B1_sel SB_T1_EAST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T1_EAST_SB_OUT_B1_sel_inst0_O)
);
SB_T1_NORTH_SB_OUT_B1_sel SB_T1_NORTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T1_NORTH_SB_OUT_B1_sel_inst0_O)
);
SB_T1_SOUTH_SB_OUT_B1_sel SB_T1_SOUTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_SOUTH_SB_OUT_B1_sel_inst0_O)
);
SB_T1_WEST_SB_OUT_B1_sel SB_T1_WEST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_WEST_SB_OUT_B1_sel_inst0_O)
);
SB_T2_EAST_SB_OUT_B1_sel SB_T2_EAST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_EAST_SB_OUT_B1_sel_inst0_O)
);
SB_T2_NORTH_SB_OUT_B1_sel SB_T2_NORTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_NORTH_SB_OUT_B1_sel_inst0_O)
);
SB_T2_SOUTH_SB_OUT_B1_sel SB_T2_SOUTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_SOUTH_SB_OUT_B1_sel_inst0_O)
);
SB_T2_WEST_SB_OUT_B1_sel SB_T2_WEST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_WEST_SB_OUT_B1_sel_inst0_O)
);
SB_T3_EAST_SB_OUT_B1_sel SB_T3_EAST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T3_EAST_SB_OUT_B1_sel_inst0_O)
);
SB_T3_NORTH_SB_OUT_B1_sel SB_T3_NORTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T3_NORTH_SB_OUT_B1_sel_inst0_O)
);
SB_T3_SOUTH_SB_OUT_B1_sel SB_T3_SOUTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T3_SOUTH_SB_OUT_B1_sel_inst0_O)
);
SB_T3_WEST_SB_OUT_B1_sel SB_T3_WEST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T3_WEST_SB_OUT_B1_sel_inst0_O)
);
SB_T4_EAST_SB_OUT_B1_sel SB_T4_EAST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T4_EAST_SB_OUT_B1_sel_inst0_O)
);
SB_T4_NORTH_SB_OUT_B1_sel SB_T4_NORTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T4_NORTH_SB_OUT_B1_sel_inst0_O)
);
SB_T4_SOUTH_SB_OUT_B1_sel SB_T4_SOUTH_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T4_SOUTH_SB_OUT_B1_sel_inst0_O)
);
SB_T4_WEST_SB_OUT_B1_sel SB_T4_WEST_SB_OUT_B1_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T4_WEST_SB_OUT_B1_sel_inst0_O)
);
MuxWrapper_1_1 WIRE_SB_T0_EAST_SB_IN_B1 (
    .I(SB_T0_EAST_SB_IN_B1),
    .O(WIRE_SB_T0_EAST_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T0_NORTH_SB_IN_B1 (
    .I(SB_T0_NORTH_SB_IN_B1),
    .O(WIRE_SB_T0_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T0_SOUTH_SB_IN_B1 (
    .I(SB_T0_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T0_WEST_SB_IN_B1 (
    .I(SB_T0_WEST_SB_IN_B1),
    .O(WIRE_SB_T0_WEST_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T1_EAST_SB_IN_B1 (
    .I(SB_T1_EAST_SB_IN_B1),
    .O(WIRE_SB_T1_EAST_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T1_NORTH_SB_IN_B1 (
    .I(SB_T1_NORTH_SB_IN_B1),
    .O(WIRE_SB_T1_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T1_SOUTH_SB_IN_B1 (
    .I(SB_T1_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T1_WEST_SB_IN_B1 (
    .I(SB_T1_WEST_SB_IN_B1),
    .O(WIRE_SB_T1_WEST_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T2_EAST_SB_IN_B1 (
    .I(SB_T2_EAST_SB_IN_B1),
    .O(WIRE_SB_T2_EAST_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T2_NORTH_SB_IN_B1 (
    .I(SB_T2_NORTH_SB_IN_B1),
    .O(WIRE_SB_T2_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T2_SOUTH_SB_IN_B1 (
    .I(SB_T2_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T2_WEST_SB_IN_B1 (
    .I(SB_T2_WEST_SB_IN_B1),
    .O(WIRE_SB_T2_WEST_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T3_EAST_SB_IN_B1 (
    .I(SB_T3_EAST_SB_IN_B1),
    .O(WIRE_SB_T3_EAST_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T3_NORTH_SB_IN_B1 (
    .I(SB_T3_NORTH_SB_IN_B1),
    .O(WIRE_SB_T3_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T3_SOUTH_SB_IN_B1 (
    .I(SB_T3_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T3_WEST_SB_IN_B1 (
    .I(SB_T3_WEST_SB_IN_B1),
    .O(WIRE_SB_T3_WEST_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T4_EAST_SB_IN_B1 (
    .I(SB_T4_EAST_SB_IN_B1),
    .O(WIRE_SB_T4_EAST_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T4_NORTH_SB_IN_B1 (
    .I(SB_T4_NORTH_SB_IN_B1),
    .O(WIRE_SB_T4_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T4_SOUTH_SB_IN_B1 (
    .I(SB_T4_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_1 WIRE_SB_T4_WEST_SB_IN_B1 (
    .I(SB_T4_WEST_SB_IN_B1),
    .O(WIRE_SB_T4_WEST_SB_IN_B1_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_28_32_inst0$bit_const_0_None (
    .out(ZextWrapper_28_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit28 ZextWrapper_28_32_inst0$self_I (
    .in(config_reg_1_O),
    .out(ZextWrapper_28_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_28_32_inst0$self_O_out;
assign ZextWrapper_28_32_inst0$self_O_out = {ZextWrapper_28_32_inst0$bit_const_0_None_out,ZextWrapper_28_32_inst0$bit_const_0_None_out,ZextWrapper_28_32_inst0$bit_const_0_None_out,ZextWrapper_28_32_inst0$bit_const_0_None_out,ZextWrapper_28_32_inst0$self_I_out[27:0]};
mantle_wire__typeBitIn32 ZextWrapper_28_32_inst0$self_O (
    .in(ZextWrapper_28_32_inst0$self_O_in),
    .out(ZextWrapper_28_32_inst0$self_O_out)
);
coreir_and #(
    .width(1)
) and1_inst0 (
    .in0(coreir_eq_1_inst0_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst0_out)
);
coreir_and #(
    .width(1)
) and1_inst1 (
    .in0(coreir_eq_1_inst1_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst1_out)
);
coreir_and #(
    .width(1)
) and1_inst10 (
    .in0(coreir_eq_1_inst10_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst10_out)
);
coreir_and #(
    .width(1)
) and1_inst11 (
    .in0(coreir_eq_1_inst11_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst11_out)
);
coreir_and #(
    .width(1)
) and1_inst12 (
    .in0(coreir_eq_1_inst12_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst12_out)
);
coreir_and #(
    .width(1)
) and1_inst13 (
    .in0(coreir_eq_1_inst13_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst13_out)
);
coreir_and #(
    .width(1)
) and1_inst14 (
    .in0(coreir_eq_1_inst14_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst14_out)
);
coreir_and #(
    .width(1)
) and1_inst15 (
    .in0(coreir_eq_1_inst15_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst15_out)
);
coreir_and #(
    .width(1)
) and1_inst16 (
    .in0(coreir_eq_1_inst16_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst16_out)
);
coreir_and #(
    .width(1)
) and1_inst17 (
    .in0(coreir_eq_1_inst17_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst17_out)
);
coreir_and #(
    .width(1)
) and1_inst18 (
    .in0(coreir_eq_1_inst18_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst18_out)
);
coreir_and #(
    .width(1)
) and1_inst19 (
    .in0(coreir_eq_1_inst19_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst19_out)
);
coreir_and #(
    .width(1)
) and1_inst2 (
    .in0(coreir_eq_1_inst2_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst2_out)
);
coreir_and #(
    .width(1)
) and1_inst3 (
    .in0(coreir_eq_1_inst3_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst3_out)
);
coreir_and #(
    .width(1)
) and1_inst4 (
    .in0(coreir_eq_1_inst4_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst4_out)
);
coreir_and #(
    .width(1)
) and1_inst5 (
    .in0(coreir_eq_1_inst5_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst5_out)
);
coreir_and #(
    .width(1)
) and1_inst6 (
    .in0(coreir_eq_1_inst6_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst6_out)
);
coreir_and #(
    .width(1)
) and1_inst7 (
    .in0(coreir_eq_1_inst7_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst7_out)
);
coreir_and #(
    .width(1)
) and1_inst8 (
    .in0(coreir_eq_1_inst8_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst8_out)
);
coreir_and #(
    .width(1)
) and1_inst9 (
    .in0(coreir_eq_1_inst9_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst9_out)
);
ConfigRegister_32_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_28_8_32_1 config_reg_1 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_1_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
coreir_const #(
    .value(1'h1),
    .width(1)
) const_1_1 (
    .out(const_1_1_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst0 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_NORTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst0_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst1 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_SOUTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst1_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst10 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_EAST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst10_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst11 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_WEST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst11_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst12 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_NORTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst12_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst13 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_SOUTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst13_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst14 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_EAST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst14_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst15 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_WEST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst15_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst16 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_NORTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst16_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst17 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_SOUTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst17_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst18 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_EAST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst18_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst19 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_WEST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst19_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst2 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_EAST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst2_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst3 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_WEST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst3_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst4 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_NORTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst4_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst5 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_SOUTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst5_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst6 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_EAST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst6_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst7 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_WEST_B1_sel_inst0_O),
    .out(coreir_eq_1_inst7_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst8 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_NORTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst8_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst9 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_SOUTH_B1_sel_inst0_O),
    .out(coreir_eq_1_inst9_out)
);
assign SB_T0_EAST_SB_OUT_B1 = RMUX_T0_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T0_NORTH_SB_OUT_B1 = RMUX_T0_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T0_SOUTH_SB_OUT_B1 = RMUX_T0_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T0_WEST_SB_OUT_B1 = RMUX_T0_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T1_EAST_SB_OUT_B1 = RMUX_T1_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T1_NORTH_SB_OUT_B1 = RMUX_T1_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T1_SOUTH_SB_OUT_B1 = RMUX_T1_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T1_WEST_SB_OUT_B1 = RMUX_T1_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T2_EAST_SB_OUT_B1 = RMUX_T2_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T2_NORTH_SB_OUT_B1 = RMUX_T2_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T2_SOUTH_SB_OUT_B1 = RMUX_T2_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T2_WEST_SB_OUT_B1 = RMUX_T2_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T3_EAST_SB_OUT_B1 = RMUX_T3_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T3_NORTH_SB_OUT_B1 = RMUX_T3_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T3_SOUTH_SB_OUT_B1 = RMUX_T3_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T3_WEST_SB_OUT_B1 = RMUX_T3_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T4_EAST_SB_OUT_B1 = RMUX_T4_EAST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T4_NORTH_SB_OUT_B1 = RMUX_T4_NORTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T4_SOUTH_SB_OUT_B1 = RMUX_T4_SOUTH_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign SB_T4_WEST_SB_OUT_B1 = RMUX_T4_WEST_B1$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
assign read_config_data = MuxWrapper_2_32_inst0$Mux2x32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
endmodule

module SB_ID0_5TRACKS_B16_PE (
    input [15:0] SB_T0_EAST_SB_IN_B16,
    output [15:0] SB_T0_EAST_SB_OUT_B16,
    input [15:0] SB_T0_NORTH_SB_IN_B16,
    output [15:0] SB_T0_NORTH_SB_OUT_B16,
    input [15:0] SB_T0_SOUTH_SB_IN_B16,
    output [15:0] SB_T0_SOUTH_SB_OUT_B16,
    input [15:0] SB_T0_WEST_SB_IN_B16,
    output [15:0] SB_T0_WEST_SB_OUT_B16,
    input [15:0] SB_T1_EAST_SB_IN_B16,
    output [15:0] SB_T1_EAST_SB_OUT_B16,
    input [15:0] SB_T1_NORTH_SB_IN_B16,
    output [15:0] SB_T1_NORTH_SB_OUT_B16,
    input [15:0] SB_T1_SOUTH_SB_IN_B16,
    output [15:0] SB_T1_SOUTH_SB_OUT_B16,
    input [15:0] SB_T1_WEST_SB_IN_B16,
    output [15:0] SB_T1_WEST_SB_OUT_B16,
    input [15:0] SB_T2_EAST_SB_IN_B16,
    output [15:0] SB_T2_EAST_SB_OUT_B16,
    input [15:0] SB_T2_NORTH_SB_IN_B16,
    output [15:0] SB_T2_NORTH_SB_OUT_B16,
    input [15:0] SB_T2_SOUTH_SB_IN_B16,
    output [15:0] SB_T2_SOUTH_SB_OUT_B16,
    input [15:0] SB_T2_WEST_SB_IN_B16,
    output [15:0] SB_T2_WEST_SB_OUT_B16,
    input [15:0] SB_T3_EAST_SB_IN_B16,
    output [15:0] SB_T3_EAST_SB_OUT_B16,
    input [15:0] SB_T3_NORTH_SB_IN_B16,
    output [15:0] SB_T3_NORTH_SB_OUT_B16,
    input [15:0] SB_T3_SOUTH_SB_IN_B16,
    output [15:0] SB_T3_SOUTH_SB_OUT_B16,
    input [15:0] SB_T3_WEST_SB_IN_B16,
    output [15:0] SB_T3_WEST_SB_OUT_B16,
    input [15:0] SB_T4_EAST_SB_IN_B16,
    output [15:0] SB_T4_EAST_SB_OUT_B16,
    input [15:0] SB_T4_NORTH_SB_IN_B16,
    output [15:0] SB_T4_NORTH_SB_OUT_B16,
    input [15:0] SB_T4_SOUTH_SB_IN_B16,
    output [15:0] SB_T4_SOUTH_SB_OUT_B16,
    input [15:0] SB_T4_WEST_SB_IN_B16,
    output [15:0] SB_T4_WEST_SB_OUT_B16,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    input [15:0] pe_outputs_0,
    output [31:0] read_config_data,
    input reset,
    input [0:0] stall
);
wire [0:0] Invert1_inst0_out;
wire [15:0] MUX_SB_T0_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out;
wire [15:0] MUX_SB_T0_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out;
wire [15:0] MUX_SB_T0_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out;
wire [15:0] MUX_SB_T0_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out;
wire [15:0] MUX_SB_T1_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out;
wire [15:0] MUX_SB_T1_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out;
wire [15:0] MUX_SB_T1_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out;
wire [15:0] MUX_SB_T1_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out;
wire [15:0] MUX_SB_T2_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out;
wire [15:0] MUX_SB_T2_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out;
wire [15:0] MUX_SB_T2_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out;
wire [15:0] MUX_SB_T2_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out;
wire [15:0] MUX_SB_T3_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out;
wire [15:0] MUX_SB_T3_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out;
wire [15:0] MUX_SB_T3_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out;
wire [15:0] MUX_SB_T3_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out;
wire [15:0] MUX_SB_T4_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out;
wire [15:0] MUX_SB_T4_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out;
wire [15:0] MUX_SB_T4_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out;
wire [15:0] MUX_SB_T4_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out;
wire [31:0] MuxWrapper_2_32_inst0$Mux2x32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
wire [15:0] REG_T0_EAST_B16_O;
wire [15:0] REG_T0_NORTH_B16_O;
wire [15:0] REG_T0_SOUTH_B16_O;
wire [15:0] REG_T0_WEST_B16_O;
wire [15:0] REG_T1_EAST_B16_O;
wire [15:0] REG_T1_NORTH_B16_O;
wire [15:0] REG_T1_SOUTH_B16_O;
wire [15:0] REG_T1_WEST_B16_O;
wire [15:0] REG_T2_EAST_B16_O;
wire [15:0] REG_T2_NORTH_B16_O;
wire [15:0] REG_T2_SOUTH_B16_O;
wire [15:0] REG_T2_WEST_B16_O;
wire [15:0] REG_T3_EAST_B16_O;
wire [15:0] REG_T3_NORTH_B16_O;
wire [15:0] REG_T3_SOUTH_B16_O;
wire [15:0] REG_T3_WEST_B16_O;
wire [15:0] REG_T4_EAST_B16_O;
wire [15:0] REG_T4_NORTH_B16_O;
wire [15:0] REG_T4_SOUTH_B16_O;
wire [15:0] REG_T4_WEST_B16_O;
wire [15:0] RMUX_T0_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T0_EAST_B16_sel_inst0_O;
wire [15:0] RMUX_T0_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T0_NORTH_B16_sel_inst0_O;
wire [15:0] RMUX_T0_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T0_SOUTH_B16_sel_inst0_O;
wire [15:0] RMUX_T0_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T0_WEST_B16_sel_inst0_O;
wire [15:0] RMUX_T1_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T1_EAST_B16_sel_inst0_O;
wire [15:0] RMUX_T1_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T1_NORTH_B16_sel_inst0_O;
wire [15:0] RMUX_T1_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T1_SOUTH_B16_sel_inst0_O;
wire [15:0] RMUX_T1_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T1_WEST_B16_sel_inst0_O;
wire [15:0] RMUX_T2_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T2_EAST_B16_sel_inst0_O;
wire [15:0] RMUX_T2_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T2_NORTH_B16_sel_inst0_O;
wire [15:0] RMUX_T2_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T2_SOUTH_B16_sel_inst0_O;
wire [15:0] RMUX_T2_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T2_WEST_B16_sel_inst0_O;
wire [15:0] RMUX_T3_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T3_EAST_B16_sel_inst0_O;
wire [15:0] RMUX_T3_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T3_NORTH_B16_sel_inst0_O;
wire [15:0] RMUX_T3_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T3_SOUTH_B16_sel_inst0_O;
wire [15:0] RMUX_T3_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T3_WEST_B16_sel_inst0_O;
wire [15:0] RMUX_T4_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T4_EAST_B16_sel_inst0_O;
wire [15:0] RMUX_T4_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T4_NORTH_B16_sel_inst0_O;
wire [15:0] RMUX_T4_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T4_SOUTH_B16_sel_inst0_O;
wire [15:0] RMUX_T4_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T4_WEST_B16_sel_inst0_O;
wire [1:0] SB_T0_EAST_SB_OUT_B16_sel_inst0_O;
wire [1:0] SB_T0_NORTH_SB_OUT_B16_sel_inst0_O;
wire [1:0] SB_T0_SOUTH_SB_OUT_B16_sel_inst0_O;
wire [1:0] SB_T0_WEST_SB_OUT_B16_sel_inst0_O;
wire [1:0] SB_T1_EAST_SB_OUT_B16_sel_inst0_O;
wire [1:0] SB_T1_NORTH_SB_OUT_B16_sel_inst0_O;
wire [1:0] SB_T1_SOUTH_SB_OUT_B16_sel_inst0_O;
wire [1:0] SB_T1_WEST_SB_OUT_B16_sel_inst0_O;
wire [1:0] SB_T2_EAST_SB_OUT_B16_sel_inst0_O;
wire [1:0] SB_T2_NORTH_SB_OUT_B16_sel_inst0_O;
wire [1:0] SB_T2_SOUTH_SB_OUT_B16_sel_inst0_O;
wire [1:0] SB_T2_WEST_SB_OUT_B16_sel_inst0_O;
wire [1:0] SB_T3_EAST_SB_OUT_B16_sel_inst0_O;
wire [1:0] SB_T3_NORTH_SB_OUT_B16_sel_inst0_O;
wire [1:0] SB_T3_SOUTH_SB_OUT_B16_sel_inst0_O;
wire [1:0] SB_T3_WEST_SB_OUT_B16_sel_inst0_O;
wire [1:0] SB_T4_EAST_SB_OUT_B16_sel_inst0_O;
wire [1:0] SB_T4_NORTH_SB_OUT_B16_sel_inst0_O;
wire [1:0] SB_T4_SOUTH_SB_OUT_B16_sel_inst0_O;
wire [1:0] SB_T4_WEST_SB_OUT_B16_sel_inst0_O;
wire [15:0] WIRE_SB_T0_EAST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T0_NORTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T0_SOUTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T0_WEST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T1_EAST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T1_NORTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T1_SOUTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T1_WEST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T2_EAST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T2_NORTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T2_SOUTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T2_WEST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T3_EAST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T3_NORTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T3_SOUTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T3_WEST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T4_EAST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T4_NORTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T4_SOUTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T4_WEST_SB_IN_B16_O;
wire ZextWrapper_28_32_inst0$bit_const_0_None_out;
wire [27:0] ZextWrapper_28_32_inst0$self_I_out;
wire [31:0] ZextWrapper_28_32_inst0$self_O_in;
wire [0:0] and1_inst0_out;
wire [0:0] and1_inst1_out;
wire [0:0] and1_inst10_out;
wire [0:0] and1_inst11_out;
wire [0:0] and1_inst12_out;
wire [0:0] and1_inst13_out;
wire [0:0] and1_inst14_out;
wire [0:0] and1_inst15_out;
wire [0:0] and1_inst16_out;
wire [0:0] and1_inst17_out;
wire [0:0] and1_inst18_out;
wire [0:0] and1_inst19_out;
wire [0:0] and1_inst2_out;
wire [0:0] and1_inst3_out;
wire [0:0] and1_inst4_out;
wire [0:0] and1_inst5_out;
wire [0:0] and1_inst6_out;
wire [0:0] and1_inst7_out;
wire [0:0] and1_inst8_out;
wire [0:0] and1_inst9_out;
wire [31:0] config_reg_0_O;
wire [27:0] config_reg_1_O;
wire [0:0] const_1_1_out;
wire coreir_eq_1_inst0_out;
wire coreir_eq_1_inst1_out;
wire coreir_eq_1_inst10_out;
wire coreir_eq_1_inst11_out;
wire coreir_eq_1_inst12_out;
wire coreir_eq_1_inst13_out;
wire coreir_eq_1_inst14_out;
wire coreir_eq_1_inst15_out;
wire coreir_eq_1_inst16_out;
wire coreir_eq_1_inst17_out;
wire coreir_eq_1_inst18_out;
wire coreir_eq_1_inst19_out;
wire coreir_eq_1_inst2_out;
wire coreir_eq_1_inst3_out;
wire coreir_eq_1_inst4_out;
wire coreir_eq_1_inst5_out;
wire coreir_eq_1_inst6_out;
wire coreir_eq_1_inst7_out;
wire coreir_eq_1_inst8_out;
wire coreir_eq_1_inst9_out;
coreir_not #(
    .width(1)
) Invert1_inst0 (
    .in(stall),
    .out(Invert1_inst0_out)
);
commonlib_muxn__N4__width16 MUX_SB_T0_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0 (
    .in_data_0(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .in_data_3(pe_outputs_0),
    .in_sel(SB_T0_EAST_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T0_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out)
);
commonlib_muxn__N4__width16 MUX_SB_T0_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0 (
    .in_data_0(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .in_data_3(pe_outputs_0),
    .in_sel(SB_T0_NORTH_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T0_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out)
);
commonlib_muxn__N4__width16 MUX_SB_T0_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0 (
    .in_data_0(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .in_data_3(pe_outputs_0),
    .in_sel(SB_T0_SOUTH_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T0_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out)
);
commonlib_muxn__N4__width16 MUX_SB_T0_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0 (
    .in_data_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .in_data_3(pe_outputs_0),
    .in_sel(SB_T0_WEST_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T0_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out)
);
commonlib_muxn__N4__width16 MUX_SB_T1_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0 (
    .in_data_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .in_data_3(pe_outputs_0),
    .in_sel(SB_T1_EAST_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T1_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out)
);
commonlib_muxn__N4__width16 MUX_SB_T1_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0 (
    .in_data_0(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .in_data_3(pe_outputs_0),
    .in_sel(SB_T1_NORTH_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T1_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out)
);
commonlib_muxn__N4__width16 MUX_SB_T1_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0 (
    .in_data_0(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .in_data_3(pe_outputs_0),
    .in_sel(SB_T1_SOUTH_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T1_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out)
);
commonlib_muxn__N4__width16 MUX_SB_T1_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0 (
    .in_data_0(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .in_data_3(pe_outputs_0),
    .in_sel(SB_T1_WEST_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T1_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out)
);
commonlib_muxn__N4__width16 MUX_SB_T2_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0 (
    .in_data_0(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .in_data_3(pe_outputs_0),
    .in_sel(SB_T2_EAST_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T2_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out)
);
commonlib_muxn__N4__width16 MUX_SB_T2_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0 (
    .in_data_0(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .in_data_3(pe_outputs_0),
    .in_sel(SB_T2_NORTH_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T2_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out)
);
commonlib_muxn__N4__width16 MUX_SB_T2_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0 (
    .in_data_0(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .in_data_3(pe_outputs_0),
    .in_sel(SB_T2_SOUTH_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T2_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out)
);
commonlib_muxn__N4__width16 MUX_SB_T2_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0 (
    .in_data_0(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .in_data_3(pe_outputs_0),
    .in_sel(SB_T2_WEST_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T2_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out)
);
commonlib_muxn__N4__width16 MUX_SB_T3_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0 (
    .in_data_0(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .in_data_3(pe_outputs_0),
    .in_sel(SB_T3_EAST_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T3_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out)
);
commonlib_muxn__N4__width16 MUX_SB_T3_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0 (
    .in_data_0(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .in_data_3(pe_outputs_0),
    .in_sel(SB_T3_NORTH_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T3_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out)
);
commonlib_muxn__N4__width16 MUX_SB_T3_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0 (
    .in_data_0(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .in_data_3(pe_outputs_0),
    .in_sel(SB_T3_SOUTH_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T3_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out)
);
commonlib_muxn__N4__width16 MUX_SB_T3_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0 (
    .in_data_0(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .in_data_3(pe_outputs_0),
    .in_sel(SB_T3_WEST_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T3_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out)
);
commonlib_muxn__N4__width16 MUX_SB_T4_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0 (
    .in_data_0(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .in_data_3(pe_outputs_0),
    .in_sel(SB_T4_EAST_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T4_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out)
);
commonlib_muxn__N4__width16 MUX_SB_T4_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0 (
    .in_data_0(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .in_data_3(pe_outputs_0),
    .in_sel(SB_T4_NORTH_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T4_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out)
);
commonlib_muxn__N4__width16 MUX_SB_T4_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0 (
    .in_data_0(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .in_data_3(pe_outputs_0),
    .in_sel(SB_T4_SOUTH_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T4_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out)
);
commonlib_muxn__N4__width16 MUX_SB_T4_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0 (
    .in_data_0(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .in_data_3(pe_outputs_0),
    .in_sel(SB_T4_WEST_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T4_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out)
);
coreir_mux #(
    .width(32)
) MuxWrapper_2_32_inst0$Mux2x32_inst0$coreir_commonlib_mux2x32_inst0$_join (
    .in0(config_reg_0_O),
    .in1(ZextWrapper_28_32_inst0$self_O_in),
    .sel(config_config_addr[0]),
    .out(MuxWrapper_2_32_inst0$Mux2x32_inst0$coreir_commonlib_mux2x32_inst0$_join_out)
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T0_EAST_B16 (
    .I(MUX_SB_T0_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .O(REG_T0_EAST_B16_O),
    .CLK(clk),
    .CE(and1_inst2_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T0_NORTH_B16 (
    .I(MUX_SB_T0_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .O(REG_T0_NORTH_B16_O),
    .CLK(clk),
    .CE(and1_inst0_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T0_SOUTH_B16 (
    .I(MUX_SB_T0_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .O(REG_T0_SOUTH_B16_O),
    .CLK(clk),
    .CE(and1_inst1_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T0_WEST_B16 (
    .I(MUX_SB_T0_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .O(REG_T0_WEST_B16_O),
    .CLK(clk),
    .CE(and1_inst3_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T1_EAST_B16 (
    .I(MUX_SB_T1_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .O(REG_T1_EAST_B16_O),
    .CLK(clk),
    .CE(and1_inst6_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T1_NORTH_B16 (
    .I(MUX_SB_T1_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .O(REG_T1_NORTH_B16_O),
    .CLK(clk),
    .CE(and1_inst4_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T1_SOUTH_B16 (
    .I(MUX_SB_T1_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .O(REG_T1_SOUTH_B16_O),
    .CLK(clk),
    .CE(and1_inst5_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T1_WEST_B16 (
    .I(MUX_SB_T1_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .O(REG_T1_WEST_B16_O),
    .CLK(clk),
    .CE(and1_inst7_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T2_EAST_B16 (
    .I(MUX_SB_T2_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .O(REG_T2_EAST_B16_O),
    .CLK(clk),
    .CE(and1_inst10_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T2_NORTH_B16 (
    .I(MUX_SB_T2_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .O(REG_T2_NORTH_B16_O),
    .CLK(clk),
    .CE(and1_inst8_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T2_SOUTH_B16 (
    .I(MUX_SB_T2_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .O(REG_T2_SOUTH_B16_O),
    .CLK(clk),
    .CE(and1_inst9_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T2_WEST_B16 (
    .I(MUX_SB_T2_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .O(REG_T2_WEST_B16_O),
    .CLK(clk),
    .CE(and1_inst11_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T3_EAST_B16 (
    .I(MUX_SB_T3_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .O(REG_T3_EAST_B16_O),
    .CLK(clk),
    .CE(and1_inst14_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T3_NORTH_B16 (
    .I(MUX_SB_T3_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .O(REG_T3_NORTH_B16_O),
    .CLK(clk),
    .CE(and1_inst12_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T3_SOUTH_B16 (
    .I(MUX_SB_T3_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .O(REG_T3_SOUTH_B16_O),
    .CLK(clk),
    .CE(and1_inst13_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T3_WEST_B16 (
    .I(MUX_SB_T3_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .O(REG_T3_WEST_B16_O),
    .CLK(clk),
    .CE(and1_inst15_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T4_EAST_B16 (
    .I(MUX_SB_T4_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .O(REG_T4_EAST_B16_O),
    .CLK(clk),
    .CE(and1_inst18_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T4_NORTH_B16 (
    .I(MUX_SB_T4_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .O(REG_T4_NORTH_B16_O),
    .CLK(clk),
    .CE(and1_inst16_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T4_SOUTH_B16 (
    .I(MUX_SB_T4_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .O(REG_T4_SOUTH_B16_O),
    .CLK(clk),
    .CE(and1_inst17_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T4_WEST_B16 (
    .I(MUX_SB_T4_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .O(REG_T4_WEST_B16_O),
    .CLK(clk),
    .CE(and1_inst19_out[0])
);
coreir_mux #(
    .width(16)
) RMUX_T0_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T0_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .in1(REG_T0_EAST_B16_O),
    .sel(RMUX_T0_EAST_B16_sel_inst0_O[0]),
    .out(RMUX_T0_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T0_EAST_B16_sel RMUX_T0_EAST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_EAST_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T0_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T0_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .in1(REG_T0_NORTH_B16_O),
    .sel(RMUX_T0_NORTH_B16_sel_inst0_O[0]),
    .out(RMUX_T0_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T0_NORTH_B16_sel RMUX_T0_NORTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_NORTH_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T0_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T0_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .in1(REG_T0_SOUTH_B16_O),
    .sel(RMUX_T0_SOUTH_B16_sel_inst0_O[0]),
    .out(RMUX_T0_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T0_SOUTH_B16_sel RMUX_T0_SOUTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_SOUTH_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T0_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T0_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .in1(REG_T0_WEST_B16_O),
    .sel(RMUX_T0_WEST_B16_sel_inst0_O[0]),
    .out(RMUX_T0_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T0_WEST_B16_sel RMUX_T0_WEST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_WEST_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T1_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T1_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .in1(REG_T1_EAST_B16_O),
    .sel(RMUX_T1_EAST_B16_sel_inst0_O[0]),
    .out(RMUX_T1_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T1_EAST_B16_sel RMUX_T1_EAST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_EAST_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T1_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T1_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .in1(REG_T1_NORTH_B16_O),
    .sel(RMUX_T1_NORTH_B16_sel_inst0_O[0]),
    .out(RMUX_T1_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T1_NORTH_B16_sel RMUX_T1_NORTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_NORTH_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T1_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T1_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .in1(REG_T1_SOUTH_B16_O),
    .sel(RMUX_T1_SOUTH_B16_sel_inst0_O[0]),
    .out(RMUX_T1_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T1_SOUTH_B16_sel RMUX_T1_SOUTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_SOUTH_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T1_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T1_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .in1(REG_T1_WEST_B16_O),
    .sel(RMUX_T1_WEST_B16_sel_inst0_O[0]),
    .out(RMUX_T1_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T1_WEST_B16_sel RMUX_T1_WEST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_WEST_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T2_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T2_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .in1(REG_T2_EAST_B16_O),
    .sel(RMUX_T2_EAST_B16_sel_inst0_O[0]),
    .out(RMUX_T2_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T2_EAST_B16_sel RMUX_T2_EAST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_EAST_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T2_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T2_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .in1(REG_T2_NORTH_B16_O),
    .sel(RMUX_T2_NORTH_B16_sel_inst0_O[0]),
    .out(RMUX_T2_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T2_NORTH_B16_sel RMUX_T2_NORTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_NORTH_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T2_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T2_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .in1(REG_T2_SOUTH_B16_O),
    .sel(RMUX_T2_SOUTH_B16_sel_inst0_O[0]),
    .out(RMUX_T2_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T2_SOUTH_B16_sel RMUX_T2_SOUTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_SOUTH_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T2_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T2_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .in1(REG_T2_WEST_B16_O),
    .sel(RMUX_T2_WEST_B16_sel_inst0_O[0]),
    .out(RMUX_T2_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T2_WEST_B16_sel RMUX_T2_WEST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_WEST_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T3_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T3_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .in1(REG_T3_EAST_B16_O),
    .sel(RMUX_T3_EAST_B16_sel_inst0_O[0]),
    .out(RMUX_T3_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T3_EAST_B16_sel RMUX_T3_EAST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_EAST_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T3_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T3_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .in1(REG_T3_NORTH_B16_O),
    .sel(RMUX_T3_NORTH_B16_sel_inst0_O[0]),
    .out(RMUX_T3_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T3_NORTH_B16_sel RMUX_T3_NORTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_NORTH_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T3_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T3_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .in1(REG_T3_SOUTH_B16_O),
    .sel(RMUX_T3_SOUTH_B16_sel_inst0_O[0]),
    .out(RMUX_T3_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T3_SOUTH_B16_sel RMUX_T3_SOUTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_SOUTH_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T3_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T3_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .in1(REG_T3_WEST_B16_O),
    .sel(RMUX_T3_WEST_B16_sel_inst0_O[0]),
    .out(RMUX_T3_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T3_WEST_B16_sel RMUX_T3_WEST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_WEST_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T4_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T4_EAST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .in1(REG_T4_EAST_B16_O),
    .sel(RMUX_T4_EAST_B16_sel_inst0_O[0]),
    .out(RMUX_T4_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T4_EAST_B16_sel RMUX_T4_EAST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_EAST_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T4_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T4_NORTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .in1(REG_T4_NORTH_B16_O),
    .sel(RMUX_T4_NORTH_B16_sel_inst0_O[0]),
    .out(RMUX_T4_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T4_NORTH_B16_sel RMUX_T4_NORTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_NORTH_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T4_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T4_SOUTH_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .in1(REG_T4_SOUTH_B16_O),
    .sel(RMUX_T4_SOUTH_B16_sel_inst0_O[0]),
    .out(RMUX_T4_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T4_SOUTH_B16_sel RMUX_T4_SOUTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_SOUTH_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T4_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T4_WEST_SB_OUT_B16$Mux4x16_inst0$coreir_commonlib_mux4x16_inst0_out),
    .in1(REG_T4_WEST_B16_O),
    .sel(RMUX_T4_WEST_B16_sel_inst0_O[0]),
    .out(RMUX_T4_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T4_WEST_B16_sel RMUX_T4_WEST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_WEST_B16_sel_inst0_O)
);
SB_T0_EAST_SB_OUT_B16_sel SB_T0_EAST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_EAST_SB_OUT_B16_sel_inst0_O)
);
SB_T0_NORTH_SB_OUT_B16_sel SB_T0_NORTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_NORTH_SB_OUT_B16_sel_inst0_O)
);
SB_T0_SOUTH_SB_OUT_B16_sel SB_T0_SOUTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_SOUTH_SB_OUT_B16_sel_inst0_O)
);
SB_T0_WEST_SB_OUT_B16_sel SB_T0_WEST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_WEST_SB_OUT_B16_sel_inst0_O)
);
SB_T1_EAST_SB_OUT_B16_sel SB_T1_EAST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T1_EAST_SB_OUT_B16_sel_inst0_O)
);
SB_T1_NORTH_SB_OUT_B16_sel SB_T1_NORTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T1_NORTH_SB_OUT_B16_sel_inst0_O)
);
SB_T1_SOUTH_SB_OUT_B16_sel SB_T1_SOUTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_SOUTH_SB_OUT_B16_sel_inst0_O)
);
SB_T1_WEST_SB_OUT_B16_sel SB_T1_WEST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_WEST_SB_OUT_B16_sel_inst0_O)
);
SB_T2_EAST_SB_OUT_B16_sel SB_T2_EAST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_EAST_SB_OUT_B16_sel_inst0_O)
);
SB_T2_NORTH_SB_OUT_B16_sel SB_T2_NORTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_NORTH_SB_OUT_B16_sel_inst0_O)
);
SB_T2_SOUTH_SB_OUT_B16_sel SB_T2_SOUTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_SOUTH_SB_OUT_B16_sel_inst0_O)
);
SB_T2_WEST_SB_OUT_B16_sel SB_T2_WEST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_WEST_SB_OUT_B16_sel_inst0_O)
);
SB_T3_EAST_SB_OUT_B16_sel SB_T3_EAST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T3_EAST_SB_OUT_B16_sel_inst0_O)
);
SB_T3_NORTH_SB_OUT_B16_sel SB_T3_NORTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T3_NORTH_SB_OUT_B16_sel_inst0_O)
);
SB_T3_SOUTH_SB_OUT_B16_sel SB_T3_SOUTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T3_SOUTH_SB_OUT_B16_sel_inst0_O)
);
SB_T3_WEST_SB_OUT_B16_sel SB_T3_WEST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T3_WEST_SB_OUT_B16_sel_inst0_O)
);
SB_T4_EAST_SB_OUT_B16_sel SB_T4_EAST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T4_EAST_SB_OUT_B16_sel_inst0_O)
);
SB_T4_NORTH_SB_OUT_B16_sel SB_T4_NORTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T4_NORTH_SB_OUT_B16_sel_inst0_O)
);
SB_T4_SOUTH_SB_OUT_B16_sel SB_T4_SOUTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T4_SOUTH_SB_OUT_B16_sel_inst0_O)
);
SB_T4_WEST_SB_OUT_B16_sel SB_T4_WEST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T4_WEST_SB_OUT_B16_sel_inst0_O)
);
MuxWrapper_1_16 WIRE_SB_T0_EAST_SB_IN_B16 (
    .I(SB_T0_EAST_SB_IN_B16),
    .O(WIRE_SB_T0_EAST_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T0_NORTH_SB_IN_B16 (
    .I(SB_T0_NORTH_SB_IN_B16),
    .O(WIRE_SB_T0_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T0_SOUTH_SB_IN_B16 (
    .I(SB_T0_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T0_WEST_SB_IN_B16 (
    .I(SB_T0_WEST_SB_IN_B16),
    .O(WIRE_SB_T0_WEST_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T1_EAST_SB_IN_B16 (
    .I(SB_T1_EAST_SB_IN_B16),
    .O(WIRE_SB_T1_EAST_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T1_NORTH_SB_IN_B16 (
    .I(SB_T1_NORTH_SB_IN_B16),
    .O(WIRE_SB_T1_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T1_SOUTH_SB_IN_B16 (
    .I(SB_T1_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T1_WEST_SB_IN_B16 (
    .I(SB_T1_WEST_SB_IN_B16),
    .O(WIRE_SB_T1_WEST_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T2_EAST_SB_IN_B16 (
    .I(SB_T2_EAST_SB_IN_B16),
    .O(WIRE_SB_T2_EAST_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T2_NORTH_SB_IN_B16 (
    .I(SB_T2_NORTH_SB_IN_B16),
    .O(WIRE_SB_T2_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T2_SOUTH_SB_IN_B16 (
    .I(SB_T2_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T2_WEST_SB_IN_B16 (
    .I(SB_T2_WEST_SB_IN_B16),
    .O(WIRE_SB_T2_WEST_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T3_EAST_SB_IN_B16 (
    .I(SB_T3_EAST_SB_IN_B16),
    .O(WIRE_SB_T3_EAST_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T3_NORTH_SB_IN_B16 (
    .I(SB_T3_NORTH_SB_IN_B16),
    .O(WIRE_SB_T3_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T3_SOUTH_SB_IN_B16 (
    .I(SB_T3_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T3_WEST_SB_IN_B16 (
    .I(SB_T3_WEST_SB_IN_B16),
    .O(WIRE_SB_T3_WEST_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T4_EAST_SB_IN_B16 (
    .I(SB_T4_EAST_SB_IN_B16),
    .O(WIRE_SB_T4_EAST_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T4_NORTH_SB_IN_B16 (
    .I(SB_T4_NORTH_SB_IN_B16),
    .O(WIRE_SB_T4_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T4_SOUTH_SB_IN_B16 (
    .I(SB_T4_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T4_WEST_SB_IN_B16 (
    .I(SB_T4_WEST_SB_IN_B16),
    .O(WIRE_SB_T4_WEST_SB_IN_B16_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_28_32_inst0$bit_const_0_None (
    .out(ZextWrapper_28_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit28 ZextWrapper_28_32_inst0$self_I (
    .in(config_reg_1_O),
    .out(ZextWrapper_28_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_28_32_inst0$self_O_out;
assign ZextWrapper_28_32_inst0$self_O_out = {ZextWrapper_28_32_inst0$bit_const_0_None_out,ZextWrapper_28_32_inst0$bit_const_0_None_out,ZextWrapper_28_32_inst0$bit_const_0_None_out,ZextWrapper_28_32_inst0$bit_const_0_None_out,ZextWrapper_28_32_inst0$self_I_out[27:0]};
mantle_wire__typeBitIn32 ZextWrapper_28_32_inst0$self_O (
    .in(ZextWrapper_28_32_inst0$self_O_in),
    .out(ZextWrapper_28_32_inst0$self_O_out)
);
coreir_and #(
    .width(1)
) and1_inst0 (
    .in0(coreir_eq_1_inst0_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst0_out)
);
coreir_and #(
    .width(1)
) and1_inst1 (
    .in0(coreir_eq_1_inst1_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst1_out)
);
coreir_and #(
    .width(1)
) and1_inst10 (
    .in0(coreir_eq_1_inst10_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst10_out)
);
coreir_and #(
    .width(1)
) and1_inst11 (
    .in0(coreir_eq_1_inst11_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst11_out)
);
coreir_and #(
    .width(1)
) and1_inst12 (
    .in0(coreir_eq_1_inst12_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst12_out)
);
coreir_and #(
    .width(1)
) and1_inst13 (
    .in0(coreir_eq_1_inst13_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst13_out)
);
coreir_and #(
    .width(1)
) and1_inst14 (
    .in0(coreir_eq_1_inst14_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst14_out)
);
coreir_and #(
    .width(1)
) and1_inst15 (
    .in0(coreir_eq_1_inst15_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst15_out)
);
coreir_and #(
    .width(1)
) and1_inst16 (
    .in0(coreir_eq_1_inst16_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst16_out)
);
coreir_and #(
    .width(1)
) and1_inst17 (
    .in0(coreir_eq_1_inst17_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst17_out)
);
coreir_and #(
    .width(1)
) and1_inst18 (
    .in0(coreir_eq_1_inst18_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst18_out)
);
coreir_and #(
    .width(1)
) and1_inst19 (
    .in0(coreir_eq_1_inst19_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst19_out)
);
coreir_and #(
    .width(1)
) and1_inst2 (
    .in0(coreir_eq_1_inst2_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst2_out)
);
coreir_and #(
    .width(1)
) and1_inst3 (
    .in0(coreir_eq_1_inst3_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst3_out)
);
coreir_and #(
    .width(1)
) and1_inst4 (
    .in0(coreir_eq_1_inst4_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst4_out)
);
coreir_and #(
    .width(1)
) and1_inst5 (
    .in0(coreir_eq_1_inst5_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst5_out)
);
coreir_and #(
    .width(1)
) and1_inst6 (
    .in0(coreir_eq_1_inst6_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst6_out)
);
coreir_and #(
    .width(1)
) and1_inst7 (
    .in0(coreir_eq_1_inst7_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst7_out)
);
coreir_and #(
    .width(1)
) and1_inst8 (
    .in0(coreir_eq_1_inst8_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst8_out)
);
coreir_and #(
    .width(1)
) and1_inst9 (
    .in0(coreir_eq_1_inst9_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst9_out)
);
ConfigRegister_32_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_28_8_32_1 config_reg_1 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_1_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
coreir_const #(
    .value(1'h1),
    .width(1)
) const_1_1 (
    .out(const_1_1_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst0 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_NORTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst0_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst1 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_SOUTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst1_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst10 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_EAST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst10_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst11 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_WEST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst11_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst12 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_NORTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst12_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst13 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_SOUTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst13_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst14 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_EAST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst14_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst15 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_WEST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst15_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst16 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_NORTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst16_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst17 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_SOUTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst17_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst18 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_EAST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst18_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst19 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_WEST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst19_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst2 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_EAST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst2_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst3 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_WEST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst3_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst4 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_NORTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst4_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst5 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_SOUTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst5_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst6 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_EAST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst6_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst7 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_WEST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst7_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst8 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_NORTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst8_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst9 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_SOUTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst9_out)
);
assign SB_T0_EAST_SB_OUT_B16 = RMUX_T0_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T0_NORTH_SB_OUT_B16 = RMUX_T0_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T0_SOUTH_SB_OUT_B16 = RMUX_T0_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T0_WEST_SB_OUT_B16 = RMUX_T0_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T1_EAST_SB_OUT_B16 = RMUX_T1_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T1_NORTH_SB_OUT_B16 = RMUX_T1_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T1_SOUTH_SB_OUT_B16 = RMUX_T1_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T1_WEST_SB_OUT_B16 = RMUX_T1_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T2_EAST_SB_OUT_B16 = RMUX_T2_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T2_NORTH_SB_OUT_B16 = RMUX_T2_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T2_SOUTH_SB_OUT_B16 = RMUX_T2_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T2_WEST_SB_OUT_B16 = RMUX_T2_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T3_EAST_SB_OUT_B16 = RMUX_T3_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T3_NORTH_SB_OUT_B16 = RMUX_T3_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T3_SOUTH_SB_OUT_B16 = RMUX_T3_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T3_WEST_SB_OUT_B16 = RMUX_T3_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T4_EAST_SB_OUT_B16 = RMUX_T4_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T4_NORTH_SB_OUT_B16 = RMUX_T4_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T4_SOUTH_SB_OUT_B16 = RMUX_T4_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T4_WEST_SB_OUT_B16 = RMUX_T4_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign read_config_data = MuxWrapper_2_32_inst0$Mux2x32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
endmodule

module ConfigRegister_27_8_32_49 (
    input clk,
    input reset,
    output [26:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [26:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0_O;
wire [7:0] const_49_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0 (
    .I(config_data[26:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h31),
    .width(8)
) const_49_8 (
    .out(const_49_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_49_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0_O;
endmodule

module ConfigRegister_27_8_32_48 (
    input clk,
    input reset,
    output [26:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [26:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0_O;
wire [7:0] const_48_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0 (
    .I(config_data[26:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h30),
    .width(8)
) const_48_8 (
    .out(const_48_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_48_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0_O;
endmodule

module ConfigRegister_27_8_32_47 (
    input clk,
    input reset,
    output [26:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [26:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0_O;
wire [7:0] const_47_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0 (
    .I(config_data[26:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h2f),
    .width(8)
) const_47_8 (
    .out(const_47_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_47_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0_O;
endmodule

module ConfigRegister_27_8_32_46 (
    input clk,
    input reset,
    output [26:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [26:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0_O;
wire [7:0] const_46_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0 (
    .I(config_data[26:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h2e),
    .width(8)
) const_46_8 (
    .out(const_46_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_46_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0_O;
endmodule

module ConfigRegister_27_8_32_45 (
    input clk,
    input reset,
    output [26:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [26:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0_O;
wire [7:0] const_45_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0 (
    .I(config_data[26:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h2d),
    .width(8)
) const_45_8 (
    .out(const_45_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_45_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0_O;
endmodule

module ConfigRegister_27_8_32_44 (
    input clk,
    input reset,
    output [26:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [26:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0_O;
wire [7:0] const_44_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0 (
    .I(config_data[26:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h2c),
    .width(8)
) const_44_8 (
    .out(const_44_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_44_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0_O;
endmodule

module ConfigRegister_27_8_32_43 (
    input clk,
    input reset,
    output [26:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [26:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0_O;
wire [7:0] const_43_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0 (
    .I(config_data[26:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h2b),
    .width(8)
) const_43_8 (
    .out(const_43_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_43_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0_O;
endmodule

module ConfigRegister_27_8_32_42 (
    input clk,
    input reset,
    output [26:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [26:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0_O;
wire [7:0] const_42_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0 (
    .I(config_data[26:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h2a),
    .width(8)
) const_42_8 (
    .out(const_42_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_42_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_27_inst0_O;
endmodule

module ConfigRegister_25_8_32_74 (
    input clk,
    input reset,
    output [24:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [24:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_25_inst0_O;
wire [7:0] const_74_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_25 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_25_inst0 (
    .I(config_data[24:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_25_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h4a),
    .width(8)
) const_74_8 (
    .out(const_74_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_74_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_25_inst0_O;
endmodule

module ConfigRegister_25_8_32_41 (
    input clk,
    input reset,
    output [24:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [24:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_25_inst0_O;
wire [7:0] const_41_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_25 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_25_inst0 (
    .I(config_data[24:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_25_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h29),
    .width(8)
) const_41_8 (
    .out(const_41_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_41_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_25_inst0_O;
endmodule

module ConfigRegister_23_8_32_4 (
    input clk,
    input reset,
    output [22:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [22:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_23_inst0_O;
wire [7:0] const_4_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_23 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_23_inst0 (
    .I(config_data[22:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_23_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h04),
    .width(8)
) const_4_8 (
    .out(const_4_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_4_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_23_inst0_O;
endmodule

module ConfigRegister_23_8_32_0 (
    input clk,
    input reset,
    output [22:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [22:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_23_inst0_O;
wire [7:0] const_0_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_23 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_23_inst0 (
    .I(config_data[22:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_23_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_0_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_23_inst0_O;
endmodule

module ConfigRegister_20_8_32_69 (
    input clk,
    input reset,
    output [19:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [19:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0_O;
wire [7:0] const_69_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0 (
    .I(config_data[19:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h45),
    .width(8)
) const_69_8 (
    .out(const_69_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_69_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0_O;
endmodule

module ConfigRegister_20_8_32_65 (
    input clk,
    input reset,
    output [19:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [19:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0_O;
wire [7:0] const_65_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0 (
    .I(config_data[19:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h41),
    .width(8)
) const_65_8 (
    .out(const_65_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_65_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0_O;
endmodule

module ConfigRegister_20_8_32_54 (
    input clk,
    input reset,
    output [19:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [19:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0_O;
wire [7:0] const_54_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0 (
    .I(config_data[19:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h36),
    .width(8)
) const_54_8 (
    .out(const_54_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_54_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0_O;
endmodule

module ConfigRegister_20_8_32_38 (
    input clk,
    input reset,
    output [19:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [19:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0_O;
wire [7:0] const_38_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0 (
    .I(config_data[19:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h26),
    .width(8)
) const_38_8 (
    .out(const_38_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_38_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0_O;
endmodule

module ConfigRegister_20_8_32_34 (
    input clk,
    input reset,
    output [19:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [19:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0_O;
wire [7:0] const_34_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0 (
    .I(config_data[19:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h22),
    .width(8)
) const_34_8 (
    .out(const_34_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_34_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0_O;
endmodule

module ConfigRegister_20_8_32_23 (
    input clk,
    input reset,
    output [19:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [19:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0_O;
wire [7:0] const_23_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0 (
    .I(config_data[19:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h17),
    .width(8)
) const_23_8 (
    .out(const_23_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_23_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0_O;
endmodule

module ConfigRegister_20_8_32_19 (
    input clk,
    input reset,
    output [19:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [19:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0_O;
wire [7:0] const_19_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0 (
    .I(config_data[19:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h13),
    .width(8)
) const_19_8 (
    .out(const_19_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_19_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_20_inst0_O;
endmodule

module ConfigRegister_18_8_32_2 (
    input clk,
    input reset,
    output [17:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [17:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_18_inst0_O;
wire [7:0] const_2_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_18 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_18_inst0 (
    .I(config_data[17:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_18_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h02),
    .width(8)
) const_2_8 (
    .out(const_2_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_2_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_18_inst0_O;
endmodule

module SB_ID0_5TRACKS_B16_MemCore (
    input [15:0] SB_T0_EAST_SB_IN_B16,
    output [15:0] SB_T0_EAST_SB_OUT_B16,
    input [15:0] SB_T0_NORTH_SB_IN_B16,
    output [15:0] SB_T0_NORTH_SB_OUT_B16,
    input [15:0] SB_T0_SOUTH_SB_IN_B16,
    output [15:0] SB_T0_SOUTH_SB_OUT_B16,
    input [15:0] SB_T0_WEST_SB_IN_B16,
    output [15:0] SB_T0_WEST_SB_OUT_B16,
    input [15:0] SB_T1_EAST_SB_IN_B16,
    output [15:0] SB_T1_EAST_SB_OUT_B16,
    input [15:0] SB_T1_NORTH_SB_IN_B16,
    output [15:0] SB_T1_NORTH_SB_OUT_B16,
    input [15:0] SB_T1_SOUTH_SB_IN_B16,
    output [15:0] SB_T1_SOUTH_SB_OUT_B16,
    input [15:0] SB_T1_WEST_SB_IN_B16,
    output [15:0] SB_T1_WEST_SB_OUT_B16,
    input [15:0] SB_T2_EAST_SB_IN_B16,
    output [15:0] SB_T2_EAST_SB_OUT_B16,
    input [15:0] SB_T2_NORTH_SB_IN_B16,
    output [15:0] SB_T2_NORTH_SB_OUT_B16,
    input [15:0] SB_T2_SOUTH_SB_IN_B16,
    output [15:0] SB_T2_SOUTH_SB_OUT_B16,
    input [15:0] SB_T2_WEST_SB_IN_B16,
    output [15:0] SB_T2_WEST_SB_OUT_B16,
    input [15:0] SB_T3_EAST_SB_IN_B16,
    output [15:0] SB_T3_EAST_SB_OUT_B16,
    input [15:0] SB_T3_NORTH_SB_IN_B16,
    output [15:0] SB_T3_NORTH_SB_OUT_B16,
    input [15:0] SB_T3_SOUTH_SB_IN_B16,
    output [15:0] SB_T3_SOUTH_SB_OUT_B16,
    input [15:0] SB_T3_WEST_SB_IN_B16,
    output [15:0] SB_T3_WEST_SB_OUT_B16,
    input [15:0] SB_T4_EAST_SB_IN_B16,
    output [15:0] SB_T4_EAST_SB_OUT_B16,
    input [15:0] SB_T4_NORTH_SB_IN_B16,
    output [15:0] SB_T4_NORTH_SB_OUT_B16,
    input [15:0] SB_T4_SOUTH_SB_IN_B16,
    output [15:0] SB_T4_SOUTH_SB_OUT_B16,
    input [15:0] SB_T4_WEST_SB_IN_B16,
    output [15:0] SB_T4_WEST_SB_OUT_B16,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    input [15:0] data_out_0,
    input [15:0] data_out_1,
    output [31:0] read_config_data,
    input reset,
    input [0:0] stall
);
wire [0:0] Invert1_inst0_out;
wire [15:0] MUX_SB_T0_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out;
wire [15:0] MUX_SB_T0_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out;
wire [15:0] MUX_SB_T0_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out;
wire [15:0] MUX_SB_T0_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out;
wire [15:0] MUX_SB_T1_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out;
wire [15:0] MUX_SB_T1_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out;
wire [15:0] MUX_SB_T1_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out;
wire [15:0] MUX_SB_T1_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out;
wire [15:0] MUX_SB_T2_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out;
wire [15:0] MUX_SB_T2_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out;
wire [15:0] MUX_SB_T2_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out;
wire [15:0] MUX_SB_T2_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out;
wire [15:0] MUX_SB_T3_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out;
wire [15:0] MUX_SB_T3_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out;
wire [15:0] MUX_SB_T3_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out;
wire [15:0] MUX_SB_T3_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out;
wire [15:0] MUX_SB_T4_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out;
wire [15:0] MUX_SB_T4_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out;
wire [15:0] MUX_SB_T4_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out;
wire [15:0] MUX_SB_T4_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out;
wire [31:0] MuxWrapper_3_32_inst0$Mux3x32_inst0$coreir_commonlib_mux3x32_inst0_out;
wire [1:0] MuxWrapper_3_32_inst0_S_in;
wire [15:0] REG_T0_EAST_B16_O;
wire [15:0] REG_T0_NORTH_B16_O;
wire [15:0] REG_T0_SOUTH_B16_O;
wire [15:0] REG_T0_WEST_B16_O;
wire [15:0] REG_T1_EAST_B16_O;
wire [15:0] REG_T1_NORTH_B16_O;
wire [15:0] REG_T1_SOUTH_B16_O;
wire [15:0] REG_T1_WEST_B16_O;
wire [15:0] REG_T2_EAST_B16_O;
wire [15:0] REG_T2_NORTH_B16_O;
wire [15:0] REG_T2_SOUTH_B16_O;
wire [15:0] REG_T2_WEST_B16_O;
wire [15:0] REG_T3_EAST_B16_O;
wire [15:0] REG_T3_NORTH_B16_O;
wire [15:0] REG_T3_SOUTH_B16_O;
wire [15:0] REG_T3_WEST_B16_O;
wire [15:0] REG_T4_EAST_B16_O;
wire [15:0] REG_T4_NORTH_B16_O;
wire [15:0] REG_T4_SOUTH_B16_O;
wire [15:0] REG_T4_WEST_B16_O;
wire [15:0] RMUX_T0_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T0_EAST_B16_sel_inst0_O;
wire [15:0] RMUX_T0_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T0_NORTH_B16_sel_inst0_O;
wire [15:0] RMUX_T0_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T0_SOUTH_B16_sel_inst0_O;
wire [15:0] RMUX_T0_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T0_WEST_B16_sel_inst0_O;
wire [15:0] RMUX_T1_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T1_EAST_B16_sel_inst0_O;
wire [15:0] RMUX_T1_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T1_NORTH_B16_sel_inst0_O;
wire [15:0] RMUX_T1_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T1_SOUTH_B16_sel_inst0_O;
wire [15:0] RMUX_T1_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T1_WEST_B16_sel_inst0_O;
wire [15:0] RMUX_T2_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T2_EAST_B16_sel_inst0_O;
wire [15:0] RMUX_T2_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T2_NORTH_B16_sel_inst0_O;
wire [15:0] RMUX_T2_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T2_SOUTH_B16_sel_inst0_O;
wire [15:0] RMUX_T2_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T2_WEST_B16_sel_inst0_O;
wire [15:0] RMUX_T3_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T3_EAST_B16_sel_inst0_O;
wire [15:0] RMUX_T3_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T3_NORTH_B16_sel_inst0_O;
wire [15:0] RMUX_T3_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T3_SOUTH_B16_sel_inst0_O;
wire [15:0] RMUX_T3_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T3_WEST_B16_sel_inst0_O;
wire [15:0] RMUX_T4_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T4_EAST_B16_sel_inst0_O;
wire [15:0] RMUX_T4_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T4_NORTH_B16_sel_inst0_O;
wire [15:0] RMUX_T4_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T4_SOUTH_B16_sel_inst0_O;
wire [15:0] RMUX_T4_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [0:0] RMUX_T4_WEST_B16_sel_inst0_O;
wire [2:0] SB_T0_EAST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T0_NORTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T0_SOUTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T0_WEST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T1_EAST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T1_NORTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T1_SOUTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T1_WEST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T2_EAST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T2_NORTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T2_SOUTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T2_WEST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T3_EAST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T3_NORTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T3_SOUTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T3_WEST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T4_EAST_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T4_NORTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T4_SOUTH_SB_OUT_B16_sel_inst0_O;
wire [2:0] SB_T4_WEST_SB_OUT_B16_sel_inst0_O;
wire [15:0] WIRE_SB_T0_EAST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T0_NORTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T0_SOUTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T0_WEST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T1_EAST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T1_NORTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T1_SOUTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T1_WEST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T2_EAST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T2_NORTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T2_SOUTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T2_WEST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T3_EAST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T3_NORTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T3_SOUTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T3_WEST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T4_EAST_SB_IN_B16_O;
wire [15:0] WIRE_SB_T4_NORTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T4_SOUTH_SB_IN_B16_O;
wire [15:0] WIRE_SB_T4_WEST_SB_IN_B16_O;
wire ZextWrapper_18_32_inst0$bit_const_0_None_out;
wire [17:0] ZextWrapper_18_32_inst0$self_I_out;
wire [31:0] ZextWrapper_18_32_inst0$self_O_in;
wire ZextWrapper_30_32_inst0$bit_const_0_None_out;
wire [29:0] ZextWrapper_30_32_inst0$self_I_out;
wire [31:0] ZextWrapper_30_32_inst0$self_O_in;
wire [0:0] and1_inst0_out;
wire [0:0] and1_inst1_out;
wire [0:0] and1_inst10_out;
wire [0:0] and1_inst11_out;
wire [0:0] and1_inst12_out;
wire [0:0] and1_inst13_out;
wire [0:0] and1_inst14_out;
wire [0:0] and1_inst15_out;
wire [0:0] and1_inst16_out;
wire [0:0] and1_inst17_out;
wire [0:0] and1_inst18_out;
wire [0:0] and1_inst19_out;
wire [0:0] and1_inst2_out;
wire [0:0] and1_inst3_out;
wire [0:0] and1_inst4_out;
wire [0:0] and1_inst5_out;
wire [0:0] and1_inst6_out;
wire [0:0] and1_inst7_out;
wire [0:0] and1_inst8_out;
wire [0:0] and1_inst9_out;
wire [31:0] config_reg_0_O;
wire [29:0] config_reg_1_O;
wire [17:0] config_reg_2_O;
wire [0:0] const_1_1_out;
wire coreir_eq_1_inst0_out;
wire coreir_eq_1_inst1_out;
wire coreir_eq_1_inst10_out;
wire coreir_eq_1_inst11_out;
wire coreir_eq_1_inst12_out;
wire coreir_eq_1_inst13_out;
wire coreir_eq_1_inst14_out;
wire coreir_eq_1_inst15_out;
wire coreir_eq_1_inst16_out;
wire coreir_eq_1_inst17_out;
wire coreir_eq_1_inst18_out;
wire coreir_eq_1_inst19_out;
wire coreir_eq_1_inst2_out;
wire coreir_eq_1_inst3_out;
wire coreir_eq_1_inst4_out;
wire coreir_eq_1_inst5_out;
wire coreir_eq_1_inst6_out;
wire coreir_eq_1_inst7_out;
wire coreir_eq_1_inst8_out;
wire coreir_eq_1_inst9_out;
wire [7:0] self_config_config_addr_out;
coreir_not #(
    .width(1)
) Invert1_inst0 (
    .in(stall),
    .out(Invert1_inst0_out)
);
commonlib_muxn__N5__width16 MUX_SB_T0_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0 (
    .in_data_0(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .in_data_3(data_out_0),
    .in_data_4(data_out_1),
    .in_sel(SB_T0_EAST_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T0_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out)
);
commonlib_muxn__N5__width16 MUX_SB_T0_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0 (
    .in_data_0(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .in_data_3(data_out_0),
    .in_data_4(data_out_1),
    .in_sel(SB_T0_NORTH_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T0_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out)
);
commonlib_muxn__N5__width16 MUX_SB_T0_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0 (
    .in_data_0(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .in_data_3(data_out_0),
    .in_data_4(data_out_1),
    .in_sel(SB_T0_SOUTH_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T0_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out)
);
commonlib_muxn__N5__width16 MUX_SB_T0_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0 (
    .in_data_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .in_data_3(data_out_0),
    .in_data_4(data_out_1),
    .in_sel(SB_T0_WEST_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T0_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out)
);
commonlib_muxn__N5__width16 MUX_SB_T1_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0 (
    .in_data_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .in_data_3(data_out_0),
    .in_data_4(data_out_1),
    .in_sel(SB_T1_EAST_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T1_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out)
);
commonlib_muxn__N5__width16 MUX_SB_T1_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0 (
    .in_data_0(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .in_data_3(data_out_0),
    .in_data_4(data_out_1),
    .in_sel(SB_T1_NORTH_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T1_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out)
);
commonlib_muxn__N5__width16 MUX_SB_T1_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0 (
    .in_data_0(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .in_data_3(data_out_0),
    .in_data_4(data_out_1),
    .in_sel(SB_T1_SOUTH_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T1_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out)
);
commonlib_muxn__N5__width16 MUX_SB_T1_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0 (
    .in_data_0(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .in_data_3(data_out_0),
    .in_data_4(data_out_1),
    .in_sel(SB_T1_WEST_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T1_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out)
);
commonlib_muxn__N5__width16 MUX_SB_T2_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0 (
    .in_data_0(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .in_data_3(data_out_0),
    .in_data_4(data_out_1),
    .in_sel(SB_T2_EAST_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T2_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out)
);
commonlib_muxn__N5__width16 MUX_SB_T2_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0 (
    .in_data_0(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .in_data_3(data_out_0),
    .in_data_4(data_out_1),
    .in_sel(SB_T2_NORTH_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T2_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out)
);
commonlib_muxn__N5__width16 MUX_SB_T2_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0 (
    .in_data_0(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .in_data_3(data_out_0),
    .in_data_4(data_out_1),
    .in_sel(SB_T2_SOUTH_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T2_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out)
);
commonlib_muxn__N5__width16 MUX_SB_T2_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0 (
    .in_data_0(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .in_data_3(data_out_0),
    .in_data_4(data_out_1),
    .in_sel(SB_T2_WEST_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T2_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out)
);
commonlib_muxn__N5__width16 MUX_SB_T3_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0 (
    .in_data_0(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .in_data_3(data_out_0),
    .in_data_4(data_out_1),
    .in_sel(SB_T3_EAST_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T3_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out)
);
commonlib_muxn__N5__width16 MUX_SB_T3_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0 (
    .in_data_0(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .in_data_3(data_out_0),
    .in_data_4(data_out_1),
    .in_sel(SB_T3_NORTH_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T3_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out)
);
commonlib_muxn__N5__width16 MUX_SB_T3_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0 (
    .in_data_0(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .in_data_3(data_out_0),
    .in_data_4(data_out_1),
    .in_sel(SB_T3_SOUTH_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T3_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out)
);
commonlib_muxn__N5__width16 MUX_SB_T3_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0 (
    .in_data_0(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .in_data_3(data_out_0),
    .in_data_4(data_out_1),
    .in_sel(SB_T3_WEST_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T3_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out)
);
commonlib_muxn__N5__width16 MUX_SB_T4_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0 (
    .in_data_0(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .in_data_3(data_out_0),
    .in_data_4(data_out_1),
    .in_sel(SB_T4_EAST_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T4_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out)
);
commonlib_muxn__N5__width16 MUX_SB_T4_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0 (
    .in_data_0(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .in_data_3(data_out_0),
    .in_data_4(data_out_1),
    .in_sel(SB_T4_NORTH_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T4_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out)
);
commonlib_muxn__N5__width16 MUX_SB_T4_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0 (
    .in_data_0(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .in_data_3(data_out_0),
    .in_data_4(data_out_1),
    .in_sel(SB_T4_SOUTH_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T4_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out)
);
commonlib_muxn__N5__width16 MUX_SB_T4_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0 (
    .in_data_0(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .in_data_1(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .in_data_2(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .in_data_3(data_out_0),
    .in_data_4(data_out_1),
    .in_sel(SB_T4_WEST_SB_OUT_B16_sel_inst0_O),
    .out(MUX_SB_T4_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out)
);
commonlib_muxn__N3__width32 MuxWrapper_3_32_inst0$Mux3x32_inst0$coreir_commonlib_mux3x32_inst0 (
    .in_data_0(config_reg_0_O),
    .in_data_1(ZextWrapper_30_32_inst0$self_O_in),
    .in_data_2(ZextWrapper_18_32_inst0$self_O_in),
    .in_sel(MuxWrapper_3_32_inst0_S_in),
    .out(MuxWrapper_3_32_inst0$Mux3x32_inst0$coreir_commonlib_mux3x32_inst0_out)
);
mantle_wire__typeBitIn2 MuxWrapper_3_32_inst0_S (
    .in(MuxWrapper_3_32_inst0_S_in),
    .out(self_config_config_addr_out[1:0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T0_EAST_B16 (
    .I(MUX_SB_T0_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .O(REG_T0_EAST_B16_O),
    .CLK(clk),
    .CE(and1_inst2_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T0_NORTH_B16 (
    .I(MUX_SB_T0_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .O(REG_T0_NORTH_B16_O),
    .CLK(clk),
    .CE(and1_inst0_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T0_SOUTH_B16 (
    .I(MUX_SB_T0_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .O(REG_T0_SOUTH_B16_O),
    .CLK(clk),
    .CE(and1_inst1_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T0_WEST_B16 (
    .I(MUX_SB_T0_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .O(REG_T0_WEST_B16_O),
    .CLK(clk),
    .CE(and1_inst3_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T1_EAST_B16 (
    .I(MUX_SB_T1_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .O(REG_T1_EAST_B16_O),
    .CLK(clk),
    .CE(and1_inst6_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T1_NORTH_B16 (
    .I(MUX_SB_T1_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .O(REG_T1_NORTH_B16_O),
    .CLK(clk),
    .CE(and1_inst4_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T1_SOUTH_B16 (
    .I(MUX_SB_T1_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .O(REG_T1_SOUTH_B16_O),
    .CLK(clk),
    .CE(and1_inst5_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T1_WEST_B16 (
    .I(MUX_SB_T1_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .O(REG_T1_WEST_B16_O),
    .CLK(clk),
    .CE(and1_inst7_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T2_EAST_B16 (
    .I(MUX_SB_T2_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .O(REG_T2_EAST_B16_O),
    .CLK(clk),
    .CE(and1_inst10_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T2_NORTH_B16 (
    .I(MUX_SB_T2_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .O(REG_T2_NORTH_B16_O),
    .CLK(clk),
    .CE(and1_inst8_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T2_SOUTH_B16 (
    .I(MUX_SB_T2_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .O(REG_T2_SOUTH_B16_O),
    .CLK(clk),
    .CE(and1_inst9_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T2_WEST_B16 (
    .I(MUX_SB_T2_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .O(REG_T2_WEST_B16_O),
    .CLK(clk),
    .CE(and1_inst11_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T3_EAST_B16 (
    .I(MUX_SB_T3_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .O(REG_T3_EAST_B16_O),
    .CLK(clk),
    .CE(and1_inst14_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T3_NORTH_B16 (
    .I(MUX_SB_T3_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .O(REG_T3_NORTH_B16_O),
    .CLK(clk),
    .CE(and1_inst12_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T3_SOUTH_B16 (
    .I(MUX_SB_T3_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .O(REG_T3_SOUTH_B16_O),
    .CLK(clk),
    .CE(and1_inst13_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T3_WEST_B16 (
    .I(MUX_SB_T3_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .O(REG_T3_WEST_B16_O),
    .CLK(clk),
    .CE(and1_inst15_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T4_EAST_B16 (
    .I(MUX_SB_T4_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .O(REG_T4_EAST_B16_O),
    .CLK(clk),
    .CE(and1_inst18_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T4_NORTH_B16 (
    .I(MUX_SB_T4_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .O(REG_T4_NORTH_B16_O),
    .CLK(clk),
    .CE(and1_inst16_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T4_SOUTH_B16 (
    .I(MUX_SB_T4_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .O(REG_T4_SOUTH_B16_O),
    .CLK(clk),
    .CE(and1_inst17_out[0])
);
Register_has_ce_True_has_reset_False_has_async_reset_False_has_async_resetn_False_type_Bits_n_16 REG_T4_WEST_B16 (
    .I(MUX_SB_T4_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .O(REG_T4_WEST_B16_O),
    .CLK(clk),
    .CE(and1_inst19_out[0])
);
coreir_mux #(
    .width(16)
) RMUX_T0_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T0_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .in1(REG_T0_EAST_B16_O),
    .sel(RMUX_T0_EAST_B16_sel_inst0_O[0]),
    .out(RMUX_T0_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T0_EAST_B16_sel RMUX_T0_EAST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_EAST_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T0_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T0_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .in1(REG_T0_NORTH_B16_O),
    .sel(RMUX_T0_NORTH_B16_sel_inst0_O[0]),
    .out(RMUX_T0_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T0_NORTH_B16_sel RMUX_T0_NORTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_NORTH_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T0_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T0_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .in1(REG_T0_SOUTH_B16_O),
    .sel(RMUX_T0_SOUTH_B16_sel_inst0_O[0]),
    .out(RMUX_T0_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T0_SOUTH_B16_sel RMUX_T0_SOUTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_SOUTH_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T0_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T0_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .in1(REG_T0_WEST_B16_O),
    .sel(RMUX_T0_WEST_B16_sel_inst0_O[0]),
    .out(RMUX_T0_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T0_WEST_B16_sel RMUX_T0_WEST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T0_WEST_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T1_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T1_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .in1(REG_T1_EAST_B16_O),
    .sel(RMUX_T1_EAST_B16_sel_inst0_O[0]),
    .out(RMUX_T1_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T1_EAST_B16_sel RMUX_T1_EAST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_EAST_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T1_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T1_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .in1(REG_T1_NORTH_B16_O),
    .sel(RMUX_T1_NORTH_B16_sel_inst0_O[0]),
    .out(RMUX_T1_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T1_NORTH_B16_sel RMUX_T1_NORTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_NORTH_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T1_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T1_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .in1(REG_T1_SOUTH_B16_O),
    .sel(RMUX_T1_SOUTH_B16_sel_inst0_O[0]),
    .out(RMUX_T1_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T1_SOUTH_B16_sel RMUX_T1_SOUTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_SOUTH_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T1_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T1_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .in1(REG_T1_WEST_B16_O),
    .sel(RMUX_T1_WEST_B16_sel_inst0_O[0]),
    .out(RMUX_T1_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T1_WEST_B16_sel RMUX_T1_WEST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T1_WEST_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T2_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T2_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .in1(REG_T2_EAST_B16_O),
    .sel(RMUX_T2_EAST_B16_sel_inst0_O[0]),
    .out(RMUX_T2_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T2_EAST_B16_sel RMUX_T2_EAST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_EAST_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T2_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T2_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .in1(REG_T2_NORTH_B16_O),
    .sel(RMUX_T2_NORTH_B16_sel_inst0_O[0]),
    .out(RMUX_T2_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T2_NORTH_B16_sel RMUX_T2_NORTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_NORTH_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T2_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T2_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .in1(REG_T2_SOUTH_B16_O),
    .sel(RMUX_T2_SOUTH_B16_sel_inst0_O[0]),
    .out(RMUX_T2_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T2_SOUTH_B16_sel RMUX_T2_SOUTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_SOUTH_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T2_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T2_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .in1(REG_T2_WEST_B16_O),
    .sel(RMUX_T2_WEST_B16_sel_inst0_O[0]),
    .out(RMUX_T2_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T2_WEST_B16_sel RMUX_T2_WEST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T2_WEST_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T3_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T3_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .in1(REG_T3_EAST_B16_O),
    .sel(RMUX_T3_EAST_B16_sel_inst0_O[0]),
    .out(RMUX_T3_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T3_EAST_B16_sel RMUX_T3_EAST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_EAST_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T3_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T3_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .in1(REG_T3_NORTH_B16_O),
    .sel(RMUX_T3_NORTH_B16_sel_inst0_O[0]),
    .out(RMUX_T3_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T3_NORTH_B16_sel RMUX_T3_NORTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_NORTH_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T3_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T3_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .in1(REG_T3_SOUTH_B16_O),
    .sel(RMUX_T3_SOUTH_B16_sel_inst0_O[0]),
    .out(RMUX_T3_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T3_SOUTH_B16_sel RMUX_T3_SOUTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_SOUTH_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T3_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T3_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .in1(REG_T3_WEST_B16_O),
    .sel(RMUX_T3_WEST_B16_sel_inst0_O[0]),
    .out(RMUX_T3_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T3_WEST_B16_sel RMUX_T3_WEST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T3_WEST_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T4_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T4_EAST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .in1(REG_T4_EAST_B16_O),
    .sel(RMUX_T4_EAST_B16_sel_inst0_O[0]),
    .out(RMUX_T4_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T4_EAST_B16_sel RMUX_T4_EAST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_EAST_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T4_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T4_NORTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .in1(REG_T4_NORTH_B16_O),
    .sel(RMUX_T4_NORTH_B16_sel_inst0_O[0]),
    .out(RMUX_T4_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T4_NORTH_B16_sel RMUX_T4_NORTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_NORTH_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T4_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T4_SOUTH_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .in1(REG_T4_SOUTH_B16_O),
    .sel(RMUX_T4_SOUTH_B16_sel_inst0_O[0]),
    .out(RMUX_T4_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T4_SOUTH_B16_sel RMUX_T4_SOUTH_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_SOUTH_B16_sel_inst0_O)
);
coreir_mux #(
    .width(16)
) RMUX_T4_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(MUX_SB_T4_WEST_SB_OUT_B16$Mux5x16_inst0$coreir_commonlib_mux5x16_inst0_out),
    .in1(REG_T4_WEST_B16_O),
    .sel(RMUX_T4_WEST_B16_sel_inst0_O[0]),
    .out(RMUX_T4_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
RMUX_T4_WEST_B16_sel RMUX_T4_WEST_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(RMUX_T4_WEST_B16_sel_inst0_O)
);
SB_T0_EAST_SB_OUT_B16_sel_unq1 SB_T0_EAST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_EAST_SB_OUT_B16_sel_inst0_O)
);
SB_T0_NORTH_SB_OUT_B16_sel_unq1 SB_T0_NORTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_NORTH_SB_OUT_B16_sel_inst0_O)
);
SB_T0_SOUTH_SB_OUT_B16_sel_unq1 SB_T0_SOUTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_SOUTH_SB_OUT_B16_sel_inst0_O)
);
SB_T0_WEST_SB_OUT_B16_sel_unq1 SB_T0_WEST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_0_O),
    .O(SB_T0_WEST_SB_OUT_B16_sel_inst0_O)
);
SB_T1_EAST_SB_OUT_B16_sel_unq1 SB_T1_EAST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_EAST_SB_OUT_B16_sel_inst0_O)
);
SB_T1_NORTH_SB_OUT_B16_sel_unq1 SB_T1_NORTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_NORTH_SB_OUT_B16_sel_inst0_O)
);
SB_T1_SOUTH_SB_OUT_B16_sel_unq1 SB_T1_SOUTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_SOUTH_SB_OUT_B16_sel_inst0_O)
);
SB_T1_WEST_SB_OUT_B16_sel_unq1 SB_T1_WEST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T1_WEST_SB_OUT_B16_sel_inst0_O)
);
SB_T2_EAST_SB_OUT_B16_sel_unq1 SB_T2_EAST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_EAST_SB_OUT_B16_sel_inst0_O)
);
SB_T2_NORTH_SB_OUT_B16_sel_unq1 SB_T2_NORTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_NORTH_SB_OUT_B16_sel_inst0_O)
);
SB_T2_SOUTH_SB_OUT_B16_sel_unq1 SB_T2_SOUTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_SOUTH_SB_OUT_B16_sel_inst0_O)
);
SB_T2_WEST_SB_OUT_B16_sel_unq1 SB_T2_WEST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T2_WEST_SB_OUT_B16_sel_inst0_O)
);
SB_T3_EAST_SB_OUT_B16_sel_unq1 SB_T3_EAST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T3_EAST_SB_OUT_B16_sel_inst0_O)
);
SB_T3_NORTH_SB_OUT_B16_sel_unq1 SB_T3_NORTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_1_O),
    .O(SB_T3_NORTH_SB_OUT_B16_sel_inst0_O)
);
SB_T3_SOUTH_SB_OUT_B16_sel_unq1 SB_T3_SOUTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T3_SOUTH_SB_OUT_B16_sel_inst0_O)
);
SB_T3_WEST_SB_OUT_B16_sel_unq1 SB_T3_WEST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T3_WEST_SB_OUT_B16_sel_inst0_O)
);
SB_T4_EAST_SB_OUT_B16_sel_unq1 SB_T4_EAST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T4_EAST_SB_OUT_B16_sel_inst0_O)
);
SB_T4_NORTH_SB_OUT_B16_sel_unq1 SB_T4_NORTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T4_NORTH_SB_OUT_B16_sel_inst0_O)
);
SB_T4_SOUTH_SB_OUT_B16_sel_unq1 SB_T4_SOUTH_SB_OUT_B16_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T4_SOUTH_SB_OUT_B16_sel_inst0_O)
);
SB_T4_WEST_SB_OUT_B16_sel_unq1 SB_T4_WEST_SB_OUT_B16_sel_inst0 (
    .I(config_reg_2_O),
    .O(SB_T4_WEST_SB_OUT_B16_sel_inst0_O)
);
MuxWrapper_1_16 WIRE_SB_T0_EAST_SB_IN_B16 (
    .I(SB_T0_EAST_SB_IN_B16),
    .O(WIRE_SB_T0_EAST_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T0_NORTH_SB_IN_B16 (
    .I(SB_T0_NORTH_SB_IN_B16),
    .O(WIRE_SB_T0_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T0_SOUTH_SB_IN_B16 (
    .I(SB_T0_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T0_WEST_SB_IN_B16 (
    .I(SB_T0_WEST_SB_IN_B16),
    .O(WIRE_SB_T0_WEST_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T1_EAST_SB_IN_B16 (
    .I(SB_T1_EAST_SB_IN_B16),
    .O(WIRE_SB_T1_EAST_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T1_NORTH_SB_IN_B16 (
    .I(SB_T1_NORTH_SB_IN_B16),
    .O(WIRE_SB_T1_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T1_SOUTH_SB_IN_B16 (
    .I(SB_T1_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T1_WEST_SB_IN_B16 (
    .I(SB_T1_WEST_SB_IN_B16),
    .O(WIRE_SB_T1_WEST_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T2_EAST_SB_IN_B16 (
    .I(SB_T2_EAST_SB_IN_B16),
    .O(WIRE_SB_T2_EAST_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T2_NORTH_SB_IN_B16 (
    .I(SB_T2_NORTH_SB_IN_B16),
    .O(WIRE_SB_T2_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T2_SOUTH_SB_IN_B16 (
    .I(SB_T2_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T2_WEST_SB_IN_B16 (
    .I(SB_T2_WEST_SB_IN_B16),
    .O(WIRE_SB_T2_WEST_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T3_EAST_SB_IN_B16 (
    .I(SB_T3_EAST_SB_IN_B16),
    .O(WIRE_SB_T3_EAST_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T3_NORTH_SB_IN_B16 (
    .I(SB_T3_NORTH_SB_IN_B16),
    .O(WIRE_SB_T3_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T3_SOUTH_SB_IN_B16 (
    .I(SB_T3_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T3_WEST_SB_IN_B16 (
    .I(SB_T3_WEST_SB_IN_B16),
    .O(WIRE_SB_T3_WEST_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T4_EAST_SB_IN_B16 (
    .I(SB_T4_EAST_SB_IN_B16),
    .O(WIRE_SB_T4_EAST_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T4_NORTH_SB_IN_B16 (
    .I(SB_T4_NORTH_SB_IN_B16),
    .O(WIRE_SB_T4_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T4_SOUTH_SB_IN_B16 (
    .I(SB_T4_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_16 WIRE_SB_T4_WEST_SB_IN_B16 (
    .I(SB_T4_WEST_SB_IN_B16),
    .O(WIRE_SB_T4_WEST_SB_IN_B16_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_18_32_inst0$bit_const_0_None (
    .out(ZextWrapper_18_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit18 ZextWrapper_18_32_inst0$self_I (
    .in(config_reg_2_O),
    .out(ZextWrapper_18_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_18_32_inst0$self_O_out;
assign ZextWrapper_18_32_inst0$self_O_out = {ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$bit_const_0_None_out,ZextWrapper_18_32_inst0$self_I_out[17:0]};
mantle_wire__typeBitIn32 ZextWrapper_18_32_inst0$self_O (
    .in(ZextWrapper_18_32_inst0$self_O_in),
    .out(ZextWrapper_18_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_30_32_inst0$bit_const_0_None (
    .out(ZextWrapper_30_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit30 ZextWrapper_30_32_inst0$self_I (
    .in(config_reg_1_O),
    .out(ZextWrapper_30_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_30_32_inst0$self_O_out;
assign ZextWrapper_30_32_inst0$self_O_out = {ZextWrapper_30_32_inst0$bit_const_0_None_out,ZextWrapper_30_32_inst0$bit_const_0_None_out,ZextWrapper_30_32_inst0$self_I_out[29:0]};
mantle_wire__typeBitIn32 ZextWrapper_30_32_inst0$self_O (
    .in(ZextWrapper_30_32_inst0$self_O_in),
    .out(ZextWrapper_30_32_inst0$self_O_out)
);
coreir_and #(
    .width(1)
) and1_inst0 (
    .in0(coreir_eq_1_inst0_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst0_out)
);
coreir_and #(
    .width(1)
) and1_inst1 (
    .in0(coreir_eq_1_inst1_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst1_out)
);
coreir_and #(
    .width(1)
) and1_inst10 (
    .in0(coreir_eq_1_inst10_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst10_out)
);
coreir_and #(
    .width(1)
) and1_inst11 (
    .in0(coreir_eq_1_inst11_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst11_out)
);
coreir_and #(
    .width(1)
) and1_inst12 (
    .in0(coreir_eq_1_inst12_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst12_out)
);
coreir_and #(
    .width(1)
) and1_inst13 (
    .in0(coreir_eq_1_inst13_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst13_out)
);
coreir_and #(
    .width(1)
) and1_inst14 (
    .in0(coreir_eq_1_inst14_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst14_out)
);
coreir_and #(
    .width(1)
) and1_inst15 (
    .in0(coreir_eq_1_inst15_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst15_out)
);
coreir_and #(
    .width(1)
) and1_inst16 (
    .in0(coreir_eq_1_inst16_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst16_out)
);
coreir_and #(
    .width(1)
) and1_inst17 (
    .in0(coreir_eq_1_inst17_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst17_out)
);
coreir_and #(
    .width(1)
) and1_inst18 (
    .in0(coreir_eq_1_inst18_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst18_out)
);
coreir_and #(
    .width(1)
) and1_inst19 (
    .in0(coreir_eq_1_inst19_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst19_out)
);
coreir_and #(
    .width(1)
) and1_inst2 (
    .in0(coreir_eq_1_inst2_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst2_out)
);
coreir_and #(
    .width(1)
) and1_inst3 (
    .in0(coreir_eq_1_inst3_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst3_out)
);
coreir_and #(
    .width(1)
) and1_inst4 (
    .in0(coreir_eq_1_inst4_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst4_out)
);
coreir_and #(
    .width(1)
) and1_inst5 (
    .in0(coreir_eq_1_inst5_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst5_out)
);
coreir_and #(
    .width(1)
) and1_inst6 (
    .in0(coreir_eq_1_inst6_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst6_out)
);
coreir_and #(
    .width(1)
) and1_inst7 (
    .in0(coreir_eq_1_inst7_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst7_out)
);
coreir_and #(
    .width(1)
) and1_inst8 (
    .in0(coreir_eq_1_inst8_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst8_out)
);
coreir_and #(
    .width(1)
) and1_inst9 (
    .in0(coreir_eq_1_inst9_out),
    .in1(Invert1_inst0_out),
    .out(and1_inst9_out)
);
ConfigRegister_32_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_30_8_32_1 config_reg_1 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_1_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_18_8_32_2 config_reg_2 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_2_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
coreir_const #(
    .value(1'h1),
    .width(1)
) const_1_1 (
    .out(const_1_1_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst0 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_NORTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst0_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst1 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_SOUTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst1_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst10 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_EAST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst10_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst11 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_WEST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst11_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst12 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_NORTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst12_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst13 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_SOUTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst13_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst14 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_EAST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst14_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst15 (
    .in0(const_1_1_out),
    .in1(RMUX_T3_WEST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst15_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst16 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_NORTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst16_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst17 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_SOUTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst17_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst18 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_EAST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst18_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst19 (
    .in0(const_1_1_out),
    .in1(RMUX_T4_WEST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst19_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst2 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_EAST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst2_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst3 (
    .in0(const_1_1_out),
    .in1(RMUX_T0_WEST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst3_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst4 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_NORTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst4_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst5 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_SOUTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst5_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst6 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_EAST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst6_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst7 (
    .in0(const_1_1_out),
    .in1(RMUX_T1_WEST_B16_sel_inst0_O),
    .out(coreir_eq_1_inst7_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst8 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_NORTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst8_out)
);
coreir_eq #(
    .width(1)
) coreir_eq_1_inst9 (
    .in0(const_1_1_out),
    .in1(RMUX_T2_SOUTH_B16_sel_inst0_O),
    .out(coreir_eq_1_inst9_out)
);
mantle_wire__typeBit8 self_config_config_addr (
    .in(config_config_addr),
    .out(self_config_config_addr_out)
);
assign SB_T0_EAST_SB_OUT_B16 = RMUX_T0_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T0_NORTH_SB_OUT_B16 = RMUX_T0_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T0_SOUTH_SB_OUT_B16 = RMUX_T0_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T0_WEST_SB_OUT_B16 = RMUX_T0_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T1_EAST_SB_OUT_B16 = RMUX_T1_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T1_NORTH_SB_OUT_B16 = RMUX_T1_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T1_SOUTH_SB_OUT_B16 = RMUX_T1_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T1_WEST_SB_OUT_B16 = RMUX_T1_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T2_EAST_SB_OUT_B16 = RMUX_T2_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T2_NORTH_SB_OUT_B16 = RMUX_T2_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T2_SOUTH_SB_OUT_B16 = RMUX_T2_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T2_WEST_SB_OUT_B16 = RMUX_T2_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T3_EAST_SB_OUT_B16 = RMUX_T3_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T3_NORTH_SB_OUT_B16 = RMUX_T3_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T3_SOUTH_SB_OUT_B16 = RMUX_T3_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T3_WEST_SB_OUT_B16 = RMUX_T3_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T4_EAST_SB_OUT_B16 = RMUX_T4_EAST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T4_NORTH_SB_OUT_B16 = RMUX_T4_NORTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T4_SOUTH_SB_OUT_B16 = RMUX_T4_SOUTH_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign SB_T4_WEST_SB_OUT_B16 = RMUX_T4_WEST_B16$Mux2x16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign read_config_data = MuxWrapper_3_32_inst0$Mux3x32_inst0$coreir_commonlib_mux3x32_inst0_out;
endmodule

module ConfigRegister_17_8_32_78 (
    input clk,
    input reset,
    output [16:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [16:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0_O;
wire [7:0] const_78_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0 (
    .I(config_data[16:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h4e),
    .width(8)
) const_78_8 (
    .out(const_78_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_78_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0_O;
endmodule

module ConfigRegister_17_8_32_61 (
    input clk,
    input reset,
    output [16:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [16:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0_O;
wire [7:0] const_61_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0 (
    .I(config_data[16:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h3d),
    .width(8)
) const_61_8 (
    .out(const_61_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_61_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0_O;
endmodule

module ConfigRegister_17_8_32_57 (
    input clk,
    input reset,
    output [16:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [16:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0_O;
wire [7:0] const_57_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0 (
    .I(config_data[16:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h39),
    .width(8)
) const_57_8 (
    .out(const_57_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_57_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0_O;
endmodule

module ConfigRegister_17_8_32_30 (
    input clk,
    input reset,
    output [16:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [16:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0_O;
wire [7:0] const_30_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0 (
    .I(config_data[16:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h1e),
    .width(8)
) const_30_8 (
    .out(const_30_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_30_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0_O;
endmodule

module ConfigRegister_17_8_32_26 (
    input clk,
    input reset,
    output [16:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [16:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0_O;
wire [7:0] const_26_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0 (
    .I(config_data[16:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h1a),
    .width(8)
) const_26_8 (
    .out(const_26_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_26_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0_O;
endmodule

module ConfigRegister_17_8_32_15 (
    input clk,
    input reset,
    output [16:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [16:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0_O;
wire [7:0] const_15_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0 (
    .I(config_data[16:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h0f),
    .width(8)
) const_15_8 (
    .out(const_15_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_15_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0_O;
endmodule

module ConfigRegister_17_8_32_11 (
    input clk,
    input reset,
    output [16:0] O,
    input [7:0] config_addr,
    input [31:0] config_data,
    input config_en
);
wire [16:0] Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0_O;
wire [7:0] const_11_8_out;
wire magma_Bit_and_inst0_out;
wire magma_Bits_8_eq_inst0_out;
Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17 Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0 (
    .I(config_data[16:0]),
    .O(Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0_O),
    .CLK(clk),
    .CE(magma_Bit_and_inst0_out),
    .ASYNCRESET(reset)
);
coreir_const #(
    .value(8'h0b),
    .width(8)
) const_11_8 (
    .out(const_11_8_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(magma_Bits_8_eq_inst0_out),
    .in1(config_en),
    .out(magma_Bit_and_inst0_out)
);
coreir_eq #(
    .width(8)
) magma_Bits_8_eq_inst0 (
    .in0(config_addr),
    .in1(const_11_8_out),
    .out(magma_Bits_8_eq_inst0_out)
);
assign O = Register_has_ce_True_has_reset_False_has_async_reset_True_has_async_resetn_False_type_Bits_n_17_inst0_O;
endmodule

module MemCore (
    input [15:0] addr_in_0,
    input [15:0] addr_in_1,
    input [15:0] chain_data_in_0,
    input [15:0] chain_data_in_1,
    input clk,
    input [7:0] config_1_config_addr,
    input [31:0] config_1_config_data,
    input [0:0] config_1_read,
    input [0:0] config_1_write,
    input [7:0] config_2_config_addr,
    input [31:0] config_2_config_data,
    input [0:0] config_2_read,
    input [0:0] config_2_write,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input config_en_0,
    input config_en_1,
    input [0:0] config_read,
    input [0:0] config_write,
    input [15:0] data_in_0,
    input [15:0] data_in_1,
    output [15:0] data_out_0,
    output [15:0] data_out_1,
    output [0:0] empty,
    input [0:0] flush,
    output [0:0] full,
    output [31:0] read_config_data,
    output [31:0] read_config_data_1,
    output [31:0] read_config_data_2,
    input [0:0] ren_in_0,
    input [0:0] ren_in_1,
    input reset,
    output [0:0] sram_ready_out,
    input [0:0] stall,
    output [0:0] stencil_valid,
    output [0:0] valid_out_0,
    output [0:0] valid_out_1,
    input [0:0] wen_in_0,
    input [0:0] wen_in_1
);
wire [0:0] AND_CONFIG_EN_SRAM_0_out;
wire [0:0] AND_CONFIG_EN_SRAM_1_out;
wire [0:0] Invert1_inst0_out;
wire [0:0] Invert1_inst1_out;
wire [0:0] LakeTop_W_inst0_sram_ready_out;
wire [31:0] LakeTop_W_inst0_config_data_out_1;
wire [0:0] LakeTop_W_inst0_empty;
wire [15:0] LakeTop_W_inst0_data_out_1;
wire [0:0] LakeTop_W_inst0_stencil_valid;
wire [15:0] LakeTop_W_inst0_data_out_0;
wire [1:0] LakeTop_W_inst0_valid_out;
wire [0:0] LakeTop_W_inst0_full;
wire [31:0] LakeTop_W_inst0_config_data_out_0;
wire [31:0] MuxWrapper_84_32_inst0$Mux84x32_inst0$coreir_commonlib_mux84x32_inst0_out;
wire [6:0] MuxWrapper_84_32_inst0_S_in;
wire [0:0] OR_CONFIG_EN_SRAM_0_out;
wire [0:0] OR_CONFIG_EN_SRAM_1_out;
wire [0:0] OR_CONFIG_RD_SRAM_out;
wire [0:0] OR_CONFIG_WR_SRAM_out;
wire [7:0] OR_config_addr_FEATURE_O;
wire [31:0] OR_config_data_FEATURE_O;
wire ZextWrapper_17_32_inst0$bit_const_0_None_out;
wire [16:0] ZextWrapper_17_32_inst0$self_I_out;
wire [31:0] ZextWrapper_17_32_inst0$self_O_in;
wire ZextWrapper_17_32_inst1$bit_const_0_None_out;
wire [16:0] ZextWrapper_17_32_inst1$self_I_out;
wire [31:0] ZextWrapper_17_32_inst1$self_O_in;
wire ZextWrapper_17_32_inst2$bit_const_0_None_out;
wire [16:0] ZextWrapper_17_32_inst2$self_I_out;
wire [31:0] ZextWrapper_17_32_inst2$self_O_in;
wire ZextWrapper_17_32_inst3$bit_const_0_None_out;
wire [16:0] ZextWrapper_17_32_inst3$self_I_out;
wire [31:0] ZextWrapper_17_32_inst3$self_O_in;
wire ZextWrapper_17_32_inst4$bit_const_0_None_out;
wire [16:0] ZextWrapper_17_32_inst4$self_I_out;
wire [31:0] ZextWrapper_17_32_inst4$self_O_in;
wire ZextWrapper_17_32_inst5$bit_const_0_None_out;
wire [16:0] ZextWrapper_17_32_inst5$self_I_out;
wire [31:0] ZextWrapper_17_32_inst5$self_O_in;
wire ZextWrapper_17_32_inst6$bit_const_0_None_out;
wire [16:0] ZextWrapper_17_32_inst6$self_I_out;
wire [31:0] ZextWrapper_17_32_inst6$self_O_in;
wire ZextWrapper_20_32_inst0$bit_const_0_None_out;
wire [19:0] ZextWrapper_20_32_inst0$self_I_out;
wire [31:0] ZextWrapper_20_32_inst0$self_O_in;
wire ZextWrapper_20_32_inst1$bit_const_0_None_out;
wire [19:0] ZextWrapper_20_32_inst1$self_I_out;
wire [31:0] ZextWrapper_20_32_inst1$self_O_in;
wire ZextWrapper_20_32_inst2$bit_const_0_None_out;
wire [19:0] ZextWrapper_20_32_inst2$self_I_out;
wire [31:0] ZextWrapper_20_32_inst2$self_O_in;
wire ZextWrapper_20_32_inst3$bit_const_0_None_out;
wire [19:0] ZextWrapper_20_32_inst3$self_I_out;
wire [31:0] ZextWrapper_20_32_inst3$self_O_in;
wire ZextWrapper_20_32_inst4$bit_const_0_None_out;
wire [19:0] ZextWrapper_20_32_inst4$self_I_out;
wire [31:0] ZextWrapper_20_32_inst4$self_O_in;
wire ZextWrapper_20_32_inst5$bit_const_0_None_out;
wire [19:0] ZextWrapper_20_32_inst5$self_I_out;
wire [31:0] ZextWrapper_20_32_inst5$self_O_in;
wire ZextWrapper_20_32_inst6$bit_const_0_None_out;
wire [19:0] ZextWrapper_20_32_inst6$self_I_out;
wire [31:0] ZextWrapper_20_32_inst6$self_O_in;
wire ZextWrapper_23_32_inst0$bit_const_0_None_out;
wire [22:0] ZextWrapper_23_32_inst0$self_I_out;
wire [31:0] ZextWrapper_23_32_inst0$self_O_in;
wire ZextWrapper_23_32_inst1$bit_const_0_None_out;
wire [22:0] ZextWrapper_23_32_inst1$self_I_out;
wire [31:0] ZextWrapper_23_32_inst1$self_O_in;
wire ZextWrapper_25_32_inst0$bit_const_0_None_out;
wire [24:0] ZextWrapper_25_32_inst0$self_I_out;
wire [31:0] ZextWrapper_25_32_inst0$self_O_in;
wire ZextWrapper_25_32_inst1$bit_const_0_None_out;
wire [24:0] ZextWrapper_25_32_inst1$self_I_out;
wire [31:0] ZextWrapper_25_32_inst1$self_O_in;
wire ZextWrapper_27_32_inst0$bit_const_0_None_out;
wire [26:0] ZextWrapper_27_32_inst0$self_I_out;
wire [31:0] ZextWrapper_27_32_inst0$self_O_in;
wire ZextWrapper_27_32_inst1$bit_const_0_None_out;
wire [26:0] ZextWrapper_27_32_inst1$self_I_out;
wire [31:0] ZextWrapper_27_32_inst1$self_O_in;
wire ZextWrapper_27_32_inst2$bit_const_0_None_out;
wire [26:0] ZextWrapper_27_32_inst2$self_I_out;
wire [31:0] ZextWrapper_27_32_inst2$self_O_in;
wire ZextWrapper_27_32_inst3$bit_const_0_None_out;
wire [26:0] ZextWrapper_27_32_inst3$self_I_out;
wire [31:0] ZextWrapper_27_32_inst3$self_O_in;
wire ZextWrapper_27_32_inst4$bit_const_0_None_out;
wire [26:0] ZextWrapper_27_32_inst4$self_I_out;
wire [31:0] ZextWrapper_27_32_inst4$self_O_in;
wire ZextWrapper_27_32_inst5$bit_const_0_None_out;
wire [26:0] ZextWrapper_27_32_inst5$self_I_out;
wire [31:0] ZextWrapper_27_32_inst5$self_O_in;
wire ZextWrapper_27_32_inst6$bit_const_0_None_out;
wire [26:0] ZextWrapper_27_32_inst6$self_I_out;
wire [31:0] ZextWrapper_27_32_inst6$self_O_in;
wire ZextWrapper_27_32_inst7$bit_const_0_None_out;
wire [26:0] ZextWrapper_27_32_inst7$self_I_out;
wire [31:0] ZextWrapper_27_32_inst7$self_O_in;
wire ZextWrapper_29_32_inst0$bit_const_0_None_out;
wire [28:0] ZextWrapper_29_32_inst0$self_I_out;
wire [31:0] ZextWrapper_29_32_inst0$self_O_in;
wire ZextWrapper_31_32_inst0$bit_const_0_None_out;
wire [30:0] ZextWrapper_31_32_inst0$self_I_out;
wire [31:0] ZextWrapper_31_32_inst0$self_O_in;
wire [0:0] chain_chain_en_inst0_O;
wire [22:0] config_reg_0_O;
wire [31:0] config_reg_1_O;
wire [31:0] config_reg_10_O;
wire [16:0] config_reg_11_O;
wire [31:0] config_reg_12_O;
wire [31:0] config_reg_13_O;
wire [31:0] config_reg_14_O;
wire [16:0] config_reg_15_O;
wire [31:0] config_reg_16_O;
wire [31:0] config_reg_17_O;
wire [31:0] config_reg_18_O;
wire [19:0] config_reg_19_O;
wire [31:0] config_reg_2_O;
wire [31:0] config_reg_20_O;
wire [31:0] config_reg_21_O;
wire [31:0] config_reg_22_O;
wire [19:0] config_reg_23_O;
wire [31:0] config_reg_24_O;
wire [31:0] config_reg_25_O;
wire [16:0] config_reg_26_O;
wire [31:0] config_reg_27_O;
wire [31:0] config_reg_28_O;
wire [31:0] config_reg_29_O;
wire [31:0] config_reg_3_O;
wire [16:0] config_reg_30_O;
wire [31:0] config_reg_31_O;
wire [31:0] config_reg_32_O;
wire [31:0] config_reg_33_O;
wire [19:0] config_reg_34_O;
wire [31:0] config_reg_35_O;
wire [31:0] config_reg_36_O;
wire [31:0] config_reg_37_O;
wire [19:0] config_reg_38_O;
wire [31:0] config_reg_39_O;
wire [22:0] config_reg_4_O;
wire [31:0] config_reg_40_O;
wire [24:0] config_reg_41_O;
wire [26:0] config_reg_42_O;
wire [26:0] config_reg_43_O;
wire [26:0] config_reg_44_O;
wire [26:0] config_reg_45_O;
wire [26:0] config_reg_46_O;
wire [26:0] config_reg_47_O;
wire [26:0] config_reg_48_O;
wire [26:0] config_reg_49_O;
wire [31:0] config_reg_5_O;
wire [30:0] config_reg_50_O;
wire [31:0] config_reg_51_O;
wire [31:0] config_reg_52_O;
wire [31:0] config_reg_53_O;
wire [19:0] config_reg_54_O;
wire [31:0] config_reg_55_O;
wire [31:0] config_reg_56_O;
wire [16:0] config_reg_57_O;
wire [31:0] config_reg_58_O;
wire [31:0] config_reg_59_O;
wire [31:0] config_reg_6_O;
wire [31:0] config_reg_60_O;
wire [16:0] config_reg_61_O;
wire [31:0] config_reg_62_O;
wire [31:0] config_reg_63_O;
wire [31:0] config_reg_64_O;
wire [19:0] config_reg_65_O;
wire [31:0] config_reg_66_O;
wire [31:0] config_reg_67_O;
wire [31:0] config_reg_68_O;
wire [19:0] config_reg_69_O;
wire [31:0] config_reg_7_O;
wire [31:0] config_reg_70_O;
wire [31:0] config_reg_71_O;
wire [31:0] config_reg_72_O;
wire [31:0] config_reg_73_O;
wire [24:0] config_reg_74_O;
wire [31:0] config_reg_75_O;
wire [31:0] config_reg_76_O;
wire [31:0] config_reg_77_O;
wire [16:0] config_reg_78_O;
wire [31:0] config_reg_79_O;
wire [31:0] config_reg_8_O;
wire [31:0] config_reg_80_O;
wire [31:0] config_reg_81_O;
wire [31:0] config_reg_82_O;
wire [28:0] config_reg_83_O;
wire [31:0] config_reg_9_O;
wire coreir_wrapInAsyncReset_inst0_out;
wire coreir_wrapOutAsyncReset_inst0_out;
wire [15:0] fifo_ctrl_fifo_depth_inst0_O;
wire [0:0] flush_reg_sel_inst0_O;
wire [0:0] flush_reg_value_inst0_O;
wire [0:0] flush_sel$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [3:0] loops_stencil_valid_dimensionality_inst0_O;
wire [15:0] loops_stencil_valid_ranges_0_inst0_O;
wire [15:0] loops_stencil_valid_ranges_1_inst0_O;
wire [15:0] loops_stencil_valid_ranges_2_inst0_O;
wire [15:0] loops_stencil_valid_ranges_3_inst0_O;
wire [15:0] loops_stencil_valid_ranges_4_inst0_O;
wire [15:0] loops_stencil_valid_ranges_5_inst0_O;
wire [1:0] mode_inst0_O;
wire [0:0] ren_in_0_reg_sel_inst0_O;
wire [0:0] ren_in_0_reg_value_inst0_O;
wire [0:0] ren_in_0_sel$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] ren_in_1_reg_sel_inst0_O;
wire [0:0] ren_in_1_reg_value_inst0_O;
wire [0:0] ren_in_1_sel$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [7:0] self_config_config_addr_out;
wire [0:0] stencil_valid_sched_gen_enable_inst0_O;
wire [15:0] stencil_valid_sched_gen_sched_addr_gen_starting_addr_inst0_O;
wire [15:0] stencil_valid_sched_gen_sched_addr_gen_strides_0_inst0_O;
wire [15:0] stencil_valid_sched_gen_sched_addr_gen_strides_1_inst0_O;
wire [15:0] stencil_valid_sched_gen_sched_addr_gen_strides_2_inst0_O;
wire [15:0] stencil_valid_sched_gen_sched_addr_gen_strides_3_inst0_O;
wire [15:0] stencil_valid_sched_gen_sched_addr_gen_strides_4_inst0_O;
wire [15:0] stencil_valid_sched_gen_sched_addr_gen_strides_5_inst0_O;
wire [3:0] strg_ub_agg_only_agg_read_addr_gen_0_starting_addr_inst0_O;
wire [3:0] strg_ub_agg_only_agg_read_addr_gen_0_strides_0_inst0_O;
wire [3:0] strg_ub_agg_only_agg_read_addr_gen_0_strides_1_inst0_O;
wire [3:0] strg_ub_agg_only_agg_read_addr_gen_0_strides_2_inst0_O;
wire [3:0] strg_ub_agg_only_agg_read_addr_gen_0_strides_3_inst0_O;
wire [3:0] strg_ub_agg_only_agg_read_addr_gen_0_strides_4_inst0_O;
wire [3:0] strg_ub_agg_only_agg_read_addr_gen_0_strides_5_inst0_O;
wire [3:0] strg_ub_agg_only_agg_read_addr_gen_1_starting_addr_inst0_O;
wire [3:0] strg_ub_agg_only_agg_read_addr_gen_1_strides_0_inst0_O;
wire [3:0] strg_ub_agg_only_agg_read_addr_gen_1_strides_1_inst0_O;
wire [3:0] strg_ub_agg_only_agg_read_addr_gen_1_strides_2_inst0_O;
wire [3:0] strg_ub_agg_only_agg_read_addr_gen_1_strides_3_inst0_O;
wire [3:0] strg_ub_agg_only_agg_read_addr_gen_1_strides_4_inst0_O;
wire [3:0] strg_ub_agg_only_agg_read_addr_gen_1_strides_5_inst0_O;
wire [3:0] strg_ub_agg_only_agg_write_addr_gen_0_starting_addr_inst0_O;
wire [3:0] strg_ub_agg_only_agg_write_addr_gen_0_strides_0_inst0_O;
wire [3:0] strg_ub_agg_only_agg_write_addr_gen_0_strides_1_inst0_O;
wire [3:0] strg_ub_agg_only_agg_write_addr_gen_0_strides_2_inst0_O;
wire [3:0] strg_ub_agg_only_agg_write_addr_gen_0_strides_3_inst0_O;
wire [3:0] strg_ub_agg_only_agg_write_addr_gen_0_strides_4_inst0_O;
wire [3:0] strg_ub_agg_only_agg_write_addr_gen_0_strides_5_inst0_O;
wire [3:0] strg_ub_agg_only_agg_write_addr_gen_1_starting_addr_inst0_O;
wire [3:0] strg_ub_agg_only_agg_write_addr_gen_1_strides_0_inst0_O;
wire [3:0] strg_ub_agg_only_agg_write_addr_gen_1_strides_1_inst0_O;
wire [3:0] strg_ub_agg_only_agg_write_addr_gen_1_strides_2_inst0_O;
wire [3:0] strg_ub_agg_only_agg_write_addr_gen_1_strides_3_inst0_O;
wire [3:0] strg_ub_agg_only_agg_write_addr_gen_1_strides_4_inst0_O;
wire [3:0] strg_ub_agg_only_agg_write_addr_gen_1_strides_5_inst0_O;
wire [0:0] strg_ub_agg_only_agg_write_sched_gen_0_enable_inst0_O;
wire [15:0] strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr_inst0_O;
wire [15:0] strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0_inst0_O;
wire [15:0] strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1_inst0_O;
wire [15:0] strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2_inst0_O;
wire [15:0] strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3_inst0_O;
wire [15:0] strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4_inst0_O;
wire [15:0] strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5_inst0_O;
wire [0:0] strg_ub_agg_only_agg_write_sched_gen_1_enable_inst0_O;
wire [15:0] strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr_inst0_O;
wire [15:0] strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0_inst0_O;
wire [15:0] strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1_inst0_O;
wire [15:0] strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2_inst0_O;
wire [15:0] strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3_inst0_O;
wire [15:0] strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4_inst0_O;
wire [15:0] strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5_inst0_O;
wire [3:0] strg_ub_agg_only_loops_in2buf_0_dimensionality_inst0_O;
wire [15:0] strg_ub_agg_only_loops_in2buf_0_ranges_0_inst0_O;
wire [15:0] strg_ub_agg_only_loops_in2buf_0_ranges_1_inst0_O;
wire [15:0] strg_ub_agg_only_loops_in2buf_0_ranges_2_inst0_O;
wire [15:0] strg_ub_agg_only_loops_in2buf_0_ranges_3_inst0_O;
wire [15:0] strg_ub_agg_only_loops_in2buf_0_ranges_4_inst0_O;
wire [15:0] strg_ub_agg_only_loops_in2buf_0_ranges_5_inst0_O;
wire [3:0] strg_ub_agg_only_loops_in2buf_1_dimensionality_inst0_O;
wire [15:0] strg_ub_agg_only_loops_in2buf_1_ranges_0_inst0_O;
wire [15:0] strg_ub_agg_only_loops_in2buf_1_ranges_1_inst0_O;
wire [15:0] strg_ub_agg_only_loops_in2buf_1_ranges_2_inst0_O;
wire [15:0] strg_ub_agg_only_loops_in2buf_1_ranges_3_inst0_O;
wire [15:0] strg_ub_agg_only_loops_in2buf_1_ranges_4_inst0_O;
wire [15:0] strg_ub_agg_only_loops_in2buf_1_ranges_5_inst0_O;
wire [0:0] strg_ub_agg_sram_shared_agg_read_sched_gen_0_enable_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5_inst0_O;
wire [0:0] strg_ub_agg_sram_shared_agg_read_sched_gen_1_enable_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5_inst0_O;
wire [3:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5_inst0_O;
wire [3:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4_inst0_O;
wire [15:0] strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5_inst0_O;
wire [8:0] strg_ub_sram_only_input_addr_gen_0_starting_addr_inst0_O;
wire [8:0] strg_ub_sram_only_input_addr_gen_0_strides_0_inst0_O;
wire [8:0] strg_ub_sram_only_input_addr_gen_0_strides_1_inst0_O;
wire [8:0] strg_ub_sram_only_input_addr_gen_0_strides_2_inst0_O;
wire [8:0] strg_ub_sram_only_input_addr_gen_0_strides_3_inst0_O;
wire [8:0] strg_ub_sram_only_input_addr_gen_0_strides_4_inst0_O;
wire [8:0] strg_ub_sram_only_input_addr_gen_0_strides_5_inst0_O;
wire [8:0] strg_ub_sram_only_input_addr_gen_1_starting_addr_inst0_O;
wire [8:0] strg_ub_sram_only_input_addr_gen_1_strides_0_inst0_O;
wire [8:0] strg_ub_sram_only_input_addr_gen_1_strides_1_inst0_O;
wire [8:0] strg_ub_sram_only_input_addr_gen_1_strides_2_inst0_O;
wire [8:0] strg_ub_sram_only_input_addr_gen_1_strides_3_inst0_O;
wire [8:0] strg_ub_sram_only_input_addr_gen_1_strides_4_inst0_O;
wire [8:0] strg_ub_sram_only_input_addr_gen_1_strides_5_inst0_O;
wire [8:0] strg_ub_sram_only_output_addr_gen_0_starting_addr_inst0_O;
wire [8:0] strg_ub_sram_only_output_addr_gen_0_strides_0_inst0_O;
wire [8:0] strg_ub_sram_only_output_addr_gen_0_strides_1_inst0_O;
wire [8:0] strg_ub_sram_only_output_addr_gen_0_strides_2_inst0_O;
wire [8:0] strg_ub_sram_only_output_addr_gen_0_strides_3_inst0_O;
wire [8:0] strg_ub_sram_only_output_addr_gen_0_strides_4_inst0_O;
wire [8:0] strg_ub_sram_only_output_addr_gen_0_strides_5_inst0_O;
wire [8:0] strg_ub_sram_only_output_addr_gen_1_starting_addr_inst0_O;
wire [8:0] strg_ub_sram_only_output_addr_gen_1_strides_0_inst0_O;
wire [8:0] strg_ub_sram_only_output_addr_gen_1_strides_1_inst0_O;
wire [8:0] strg_ub_sram_only_output_addr_gen_1_strides_2_inst0_O;
wire [8:0] strg_ub_sram_only_output_addr_gen_1_strides_3_inst0_O;
wire [8:0] strg_ub_sram_only_output_addr_gen_1_strides_4_inst0_O;
wire [8:0] strg_ub_sram_only_output_addr_gen_1_strides_5_inst0_O;
wire [3:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5_inst0_O;
wire [3:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5_inst0_O;
wire [0:0] strg_ub_sram_tb_shared_output_sched_gen_0_enable_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5_inst0_O;
wire [0:0] strg_ub_sram_tb_shared_output_sched_gen_1_enable_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4_inst0_O;
wire [15:0] strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5_inst0_O;
wire [3:0] strg_ub_tb_only_loops_buf2out_read_0_dimensionality_inst0_O;
wire [15:0] strg_ub_tb_only_loops_buf2out_read_0_ranges_0_inst0_O;
wire [15:0] strg_ub_tb_only_loops_buf2out_read_0_ranges_1_inst0_O;
wire [15:0] strg_ub_tb_only_loops_buf2out_read_0_ranges_2_inst0_O;
wire [15:0] strg_ub_tb_only_loops_buf2out_read_0_ranges_3_inst0_O;
wire [15:0] strg_ub_tb_only_loops_buf2out_read_0_ranges_4_inst0_O;
wire [15:0] strg_ub_tb_only_loops_buf2out_read_0_ranges_5_inst0_O;
wire [3:0] strg_ub_tb_only_loops_buf2out_read_1_dimensionality_inst0_O;
wire [15:0] strg_ub_tb_only_loops_buf2out_read_1_ranges_0_inst0_O;
wire [15:0] strg_ub_tb_only_loops_buf2out_read_1_ranges_1_inst0_O;
wire [15:0] strg_ub_tb_only_loops_buf2out_read_1_ranges_2_inst0_O;
wire [15:0] strg_ub_tb_only_loops_buf2out_read_1_ranges_3_inst0_O;
wire [15:0] strg_ub_tb_only_loops_buf2out_read_1_ranges_4_inst0_O;
wire [15:0] strg_ub_tb_only_loops_buf2out_read_1_ranges_5_inst0_O;
wire [3:0] strg_ub_tb_only_tb_read_addr_gen_0_starting_addr_inst0_O;
wire [3:0] strg_ub_tb_only_tb_read_addr_gen_0_strides_0_inst0_O;
wire [3:0] strg_ub_tb_only_tb_read_addr_gen_0_strides_1_inst0_O;
wire [3:0] strg_ub_tb_only_tb_read_addr_gen_0_strides_2_inst0_O;
wire [3:0] strg_ub_tb_only_tb_read_addr_gen_0_strides_3_inst0_O;
wire [3:0] strg_ub_tb_only_tb_read_addr_gen_0_strides_4_inst0_O;
wire [3:0] strg_ub_tb_only_tb_read_addr_gen_0_strides_5_inst0_O;
wire [3:0] strg_ub_tb_only_tb_read_addr_gen_1_starting_addr_inst0_O;
wire [3:0] strg_ub_tb_only_tb_read_addr_gen_1_strides_0_inst0_O;
wire [3:0] strg_ub_tb_only_tb_read_addr_gen_1_strides_1_inst0_O;
wire [3:0] strg_ub_tb_only_tb_read_addr_gen_1_strides_2_inst0_O;
wire [3:0] strg_ub_tb_only_tb_read_addr_gen_1_strides_3_inst0_O;
wire [3:0] strg_ub_tb_only_tb_read_addr_gen_1_strides_4_inst0_O;
wire [3:0] strg_ub_tb_only_tb_read_addr_gen_1_strides_5_inst0_O;
wire [0:0] strg_ub_tb_only_tb_read_sched_gen_0_enable_inst0_O;
wire [15:0] strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr_inst0_O;
wire [15:0] strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0_inst0_O;
wire [15:0] strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1_inst0_O;
wire [15:0] strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2_inst0_O;
wire [15:0] strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3_inst0_O;
wire [15:0] strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4_inst0_O;
wire [15:0] strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5_inst0_O;
wire [0:0] strg_ub_tb_only_tb_read_sched_gen_1_enable_inst0_O;
wire [15:0] strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr_inst0_O;
wire [15:0] strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0_inst0_O;
wire [15:0] strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1_inst0_O;
wire [15:0] strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2_inst0_O;
wire [15:0] strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3_inst0_O;
wire [15:0] strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4_inst0_O;
wire [15:0] strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5_inst0_O;
wire [3:0] strg_ub_tb_only_tb_write_addr_gen_0_starting_addr_inst0_O;
wire [3:0] strg_ub_tb_only_tb_write_addr_gen_0_strides_0_inst0_O;
wire [3:0] strg_ub_tb_only_tb_write_addr_gen_0_strides_1_inst0_O;
wire [3:0] strg_ub_tb_only_tb_write_addr_gen_0_strides_2_inst0_O;
wire [3:0] strg_ub_tb_only_tb_write_addr_gen_0_strides_3_inst0_O;
wire [3:0] strg_ub_tb_only_tb_write_addr_gen_0_strides_4_inst0_O;
wire [3:0] strg_ub_tb_only_tb_write_addr_gen_0_strides_5_inst0_O;
wire [3:0] strg_ub_tb_only_tb_write_addr_gen_1_starting_addr_inst0_O;
wire [3:0] strg_ub_tb_only_tb_write_addr_gen_1_strides_0_inst0_O;
wire [3:0] strg_ub_tb_only_tb_write_addr_gen_1_strides_1_inst0_O;
wire [3:0] strg_ub_tb_only_tb_write_addr_gen_1_strides_2_inst0_O;
wire [3:0] strg_ub_tb_only_tb_write_addr_gen_1_strides_3_inst0_O;
wire [3:0] strg_ub_tb_only_tb_write_addr_gen_1_strides_4_inst0_O;
wire [3:0] strg_ub_tb_only_tb_write_addr_gen_1_strides_5_inst0_O;
wire [0:0] tile_en_inst0_O;
wire [0:0] wen_in_0_reg_sel_inst0_O;
wire [0:0] wen_in_0_reg_value_inst0_O;
wire [0:0] wen_in_0_sel$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] wen_in_1_reg_sel_inst0_O;
wire [0:0] wen_in_1_reg_value_inst0_O;
wire [0:0] wen_in_1_sel$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
coreir_and #(
    .width(1)
) AND_CONFIG_EN_SRAM_0 (
    .in0(OR_CONFIG_EN_SRAM_0_out),
    .in1(config_en_0),
    .out(AND_CONFIG_EN_SRAM_0_out)
);
coreir_and #(
    .width(1)
) AND_CONFIG_EN_SRAM_1 (
    .in0(OR_CONFIG_EN_SRAM_1_out),
    .in1(config_en_1),
    .out(AND_CONFIG_EN_SRAM_1_out)
);
coreir_not #(
    .width(1)
) Invert1_inst0 (
    .in(coreir_wrapInAsyncReset_inst0_out),
    .out(Invert1_inst0_out)
);
coreir_not #(
    .width(1)
) Invert1_inst1 (
    .in(stall),
    .out(Invert1_inst1_out)
);
wire [1:0] LakeTop_W_inst0_ren_in;
assign LakeTop_W_inst0_ren_in = {ren_in_1_sel$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0],ren_in_0_sel$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]};
wire [1:0] LakeTop_W_inst0_wen_in;
assign LakeTop_W_inst0_wen_in = {wen_in_1_sel$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0],wen_in_0_sel$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]};
wire [1:0] LakeTop_W_inst0_config_en;
assign LakeTop_W_inst0_config_en = {AND_CONFIG_EN_SRAM_1_out[0],AND_CONFIG_EN_SRAM_0_out[0]};
LakeTop_W LakeTop_W_inst0 (
    .strg_ub_agg_only_agg_write_addr_gen_0_strides_2(strg_ub_agg_only_agg_write_addr_gen_0_strides_2_inst0_O),
    .strg_ub_tb_only_loops_buf2out_read_1_dimensionality(strg_ub_tb_only_loops_buf2out_read_1_dimensionality_inst0_O),
    .strg_ub_tb_only_tb_read_addr_gen_1_starting_addr(strg_ub_tb_only_tb_read_addr_gen_1_starting_addr_inst0_O),
    .strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4(strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4_inst0_O),
    .strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1(strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1_inst0_O),
    .strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr_inst0_O),
    .strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1_inst0_O),
    .strg_ub_agg_only_agg_read_addr_gen_1_strides_1(strg_ub_agg_only_agg_read_addr_gen_1_strides_1_inst0_O),
    .strg_ub_sram_only_output_addr_gen_1_strides_3(strg_ub_sram_only_output_addr_gen_1_strides_3_inst0_O),
    .strg_ub_tb_only_tb_read_sched_gen_1_enable(strg_ub_tb_only_tb_read_sched_gen_1_enable_inst0_O),
    .addr_in_1(addr_in_1),
    .strg_ub_sram_only_input_addr_gen_1_strides_4(strg_ub_sram_only_input_addr_gen_1_strides_4_inst0_O),
    .strg_ub_sram_only_output_addr_gen_0_strides_3(strg_ub_sram_only_output_addr_gen_0_strides_3_inst0_O),
    .strg_ub_tb_only_loops_buf2out_read_0_ranges_3(strg_ub_tb_only_loops_buf2out_read_0_ranges_3_inst0_O),
    .strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4(strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4_inst0_O),
    .loops_stencil_valid_ranges_1(loops_stencil_valid_ranges_1_inst0_O),
    .strg_ub_sram_only_output_addr_gen_0_strides_5(strg_ub_sram_only_output_addr_gen_0_strides_5_inst0_O),
    .strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3(strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3_inst0_O),
    .strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2(strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2_inst0_O),
    .strg_ub_sram_only_input_addr_gen_0_strides_4(strg_ub_sram_only_input_addr_gen_0_strides_4_inst0_O),
    .strg_ub_agg_only_agg_write_addr_gen_1_strides_3(strg_ub_agg_only_agg_write_addr_gen_1_strides_3_inst0_O),
    .strg_ub_tb_only_loops_buf2out_read_1_ranges_1(strg_ub_tb_only_loops_buf2out_read_1_ranges_1_inst0_O),
    .strg_ub_tb_only_tb_write_addr_gen_0_starting_addr(strg_ub_tb_only_tb_write_addr_gen_0_starting_addr_inst0_O),
    .strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3(strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3_inst0_O),
    .strg_ub_sram_only_input_addr_gen_1_strides_3(strg_ub_sram_only_input_addr_gen_1_strides_3_inst0_O),
    .strg_ub_tb_only_tb_write_addr_gen_1_strides_3(strg_ub_tb_only_tb_write_addr_gen_1_strides_3_inst0_O),
    .strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1(strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1_inst0_O),
    .strg_ub_sram_only_output_addr_gen_1_strides_0(strg_ub_sram_only_output_addr_gen_1_strides_0_inst0_O),
    .strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4(strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4_inst0_O),
    .strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1(strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1_inst0_O),
    .chain_chain_en(chain_chain_en_inst0_O),
    .strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5_inst0_O),
    .sram_ready_out(LakeTop_W_inst0_sram_ready_out),
    .strg_ub_tb_only_tb_write_addr_gen_0_strides_0(strg_ub_tb_only_tb_write_addr_gen_0_strides_0_inst0_O),
    .tile_en(tile_en_inst0_O),
    .strg_ub_tb_only_tb_write_addr_gen_1_strides_0(strg_ub_tb_only_tb_write_addr_gen_1_strides_0_inst0_O),
    .strg_ub_sram_only_input_addr_gen_0_strides_2(strg_ub_sram_only_input_addr_gen_0_strides_2_inst0_O),
    .strg_ub_agg_only_agg_write_addr_gen_1_starting_addr(strg_ub_agg_only_agg_write_addr_gen_1_starting_addr_inst0_O),
    .strg_ub_sram_only_input_addr_gen_0_strides_5(strg_ub_sram_only_input_addr_gen_0_strides_5_inst0_O),
    .strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4(strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4_inst0_O),
    .strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0(strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0_inst0_O),
    .strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2_inst0_O),
    .strg_ub_sram_only_output_addr_gen_0_starting_addr(strg_ub_sram_only_output_addr_gen_0_starting_addr_inst0_O),
    .strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0(strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0_inst0_O),
    .strg_ub_agg_only_loops_in2buf_0_ranges_0(strg_ub_agg_only_loops_in2buf_0_ranges_0_inst0_O),
    .strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3_inst0_O),
    .strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3(strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3_inst0_O),
    .stencil_valid_sched_gen_enable(stencil_valid_sched_gen_enable_inst0_O),
    .strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality_inst0_O),
    .stencil_valid_sched_gen_sched_addr_gen_starting_addr(stencil_valid_sched_gen_sched_addr_gen_starting_addr_inst0_O),
    .strg_ub_sram_only_input_addr_gen_0_strides_3(strg_ub_sram_only_input_addr_gen_0_strides_3_inst0_O),
    .strg_ub_sram_only_output_addr_gen_1_starting_addr(strg_ub_sram_only_output_addr_gen_1_starting_addr_inst0_O),
    .strg_ub_sram_only_output_addr_gen_1_strides_4(strg_ub_sram_only_output_addr_gen_1_strides_4_inst0_O),
    .strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1_inst0_O),
    .strg_ub_sram_only_output_addr_gen_1_strides_5(strg_ub_sram_only_output_addr_gen_1_strides_5_inst0_O),
    .strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2(strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2_inst0_O),
    .strg_ub_agg_only_loops_in2buf_1_ranges_3(strg_ub_agg_only_loops_in2buf_1_ranges_3_inst0_O),
    .strg_ub_sram_only_input_addr_gen_0_strides_1(strg_ub_sram_only_input_addr_gen_0_strides_1_inst0_O),
    .stencil_valid_sched_gen_sched_addr_gen_strides_0(stencil_valid_sched_gen_sched_addr_gen_strides_0_inst0_O),
    .strg_ub_agg_only_agg_read_addr_gen_1_strides_0(strg_ub_agg_only_agg_read_addr_gen_1_strides_0_inst0_O),
    .strg_ub_agg_only_agg_read_addr_gen_0_strides_1(strg_ub_agg_only_agg_read_addr_gen_0_strides_1_inst0_O),
    .strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1(strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1_inst0_O),
    .config_data_out_1(LakeTop_W_inst0_config_data_out_1),
    .strg_ub_agg_only_loops_in2buf_0_ranges_1(strg_ub_agg_only_loops_in2buf_0_ranges_1_inst0_O),
    .strg_ub_agg_only_agg_write_addr_gen_0_strides_3(strg_ub_agg_only_agg_write_addr_gen_0_strides_3_inst0_O),
    .empty(LakeTop_W_inst0_empty),
    .strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5(strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5_inst0_O),
    .strg_ub_agg_sram_shared_agg_read_sched_gen_1_enable(strg_ub_agg_sram_shared_agg_read_sched_gen_1_enable_inst0_O),
    .strg_ub_agg_only_agg_write_addr_gen_1_strides_1(strg_ub_agg_only_agg_write_addr_gen_1_strides_1_inst0_O),
    .strg_ub_agg_only_agg_write_sched_gen_0_enable(strg_ub_agg_only_agg_write_sched_gen_0_enable_inst0_O),
    .rst_n(coreir_wrapOutAsyncReset_inst0_out),
    .strg_ub_sram_only_input_addr_gen_1_strides_0(strg_ub_sram_only_input_addr_gen_1_strides_0_inst0_O),
    .strg_ub_sram_only_input_addr_gen_1_strides_2(strg_ub_sram_only_input_addr_gen_1_strides_2_inst0_O),
    .strg_ub_tb_only_loops_buf2out_read_0_dimensionality(strg_ub_tb_only_loops_buf2out_read_0_dimensionality_inst0_O),
    .strg_ub_agg_only_loops_in2buf_0_ranges_4(strg_ub_agg_only_loops_in2buf_0_ranges_4_inst0_O),
    .strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr_inst0_O),
    .strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5(strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5_inst0_O),
    .strg_ub_sram_only_input_addr_gen_1_starting_addr(strg_ub_sram_only_input_addr_gen_1_starting_addr_inst0_O),
    .strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality_inst0_O),
    .strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5(strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5_inst0_O),
    .strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3(strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3_inst0_O),
    .strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3_inst0_O),
    .loops_stencil_valid_ranges_2(loops_stencil_valid_ranges_2_inst0_O),
    .strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2_inst0_O),
    .strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5(strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5_inst0_O),
    .clk(clk),
    .strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0_inst0_O),
    .strg_ub_tb_only_tb_write_addr_gen_0_strides_4(strg_ub_tb_only_tb_write_addr_gen_0_strides_4_inst0_O),
    .strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4(strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4_inst0_O),
    .strg_ub_sram_tb_shared_output_sched_gen_1_enable(strg_ub_sram_tb_shared_output_sched_gen_1_enable_inst0_O),
    .ren_in(LakeTop_W_inst0_ren_in),
    .strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2(strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2_inst0_O),
    .strg_ub_tb_only_tb_read_addr_gen_0_strides_5(strg_ub_tb_only_tb_read_addr_gen_0_strides_5_inst0_O),
    .data_out_1(LakeTop_W_inst0_data_out_1),
    .strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1(strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1_inst0_O),
    .data_in_1(data_in_1),
    .strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1_inst0_O),
    .strg_ub_agg_only_agg_read_addr_gen_0_strides_4(strg_ub_agg_only_agg_read_addr_gen_0_strides_4_inst0_O),
    .loops_stencil_valid_ranges_0(loops_stencil_valid_ranges_0_inst0_O),
    .strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3(strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3_inst0_O),
    .data_in_0(data_in_0),
    .mode(mode_inst0_O),
    .strg_ub_agg_only_agg_write_addr_gen_0_strides_0(strg_ub_agg_only_agg_write_addr_gen_0_strides_0_inst0_O),
    .strg_ub_agg_only_agg_write_addr_gen_1_strides_0(strg_ub_agg_only_agg_write_addr_gen_1_strides_0_inst0_O),
    .strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4(strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4_inst0_O),
    .strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5_inst0_O),
    .strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0_inst0_O),
    .strg_ub_agg_only_agg_read_addr_gen_0_strides_5(strg_ub_agg_only_agg_read_addr_gen_0_strides_5_inst0_O),
    .flush(flush_sel$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out),
    .strg_ub_agg_only_agg_write_addr_gen_0_strides_5(strg_ub_agg_only_agg_write_addr_gen_0_strides_5_inst0_O),
    .strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4_inst0_O),
    .clk_en(Invert1_inst1_out),
    .strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5_inst0_O),
    .strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2(strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2_inst0_O),
    .strg_ub_sram_only_output_addr_gen_1_strides_1(strg_ub_sram_only_output_addr_gen_1_strides_1_inst0_O),
    .strg_ub_tb_only_tb_read_sched_gen_0_enable(strg_ub_tb_only_tb_read_sched_gen_0_enable_inst0_O),
    .strg_ub_agg_only_agg_read_addr_gen_0_strides_2(strg_ub_agg_only_agg_read_addr_gen_0_strides_2_inst0_O),
    .loops_stencil_valid_ranges_4(loops_stencil_valid_ranges_4_inst0_O),
    .strg_ub_agg_only_agg_write_addr_gen_1_strides_2(strg_ub_agg_only_agg_write_addr_gen_1_strides_2_inst0_O),
    .strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2(strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2_inst0_O),
    .strg_ub_agg_only_loops_in2buf_0_ranges_3(strg_ub_agg_only_loops_in2buf_0_ranges_3_inst0_O),
    .strg_ub_sram_only_input_addr_gen_0_starting_addr(strg_ub_sram_only_input_addr_gen_0_starting_addr_inst0_O),
    .strg_ub_sram_only_input_addr_gen_1_strides_1(strg_ub_sram_only_input_addr_gen_1_strides_1_inst0_O),
    .strg_ub_tb_only_tb_write_addr_gen_0_strides_2(strg_ub_tb_only_tb_write_addr_gen_0_strides_2_inst0_O),
    .strg_ub_agg_only_loops_in2buf_1_ranges_1(strg_ub_agg_only_loops_in2buf_1_ranges_1_inst0_O),
    .strg_ub_sram_only_output_addr_gen_0_strides_2(strg_ub_sram_only_output_addr_gen_0_strides_2_inst0_O),
    .wen_in(LakeTop_W_inst0_wen_in),
    .strg_ub_agg_only_agg_write_addr_gen_0_strides_1(strg_ub_agg_only_agg_write_addr_gen_0_strides_1_inst0_O),
    .strg_ub_sram_only_input_addr_gen_1_strides_5(strg_ub_sram_only_input_addr_gen_1_strides_5_inst0_O),
    .strg_ub_agg_only_agg_read_addr_gen_0_starting_addr(strg_ub_agg_only_agg_read_addr_gen_0_starting_addr_inst0_O),
    .strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4_inst0_O),
    .strg_ub_agg_only_agg_read_addr_gen_1_strides_2(strg_ub_agg_only_agg_read_addr_gen_1_strides_2_inst0_O),
    .strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1(strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1_inst0_O),
    .strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1(strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1_inst0_O),
    .loops_stencil_valid_ranges_3(loops_stencil_valid_ranges_3_inst0_O),
    .strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2_inst0_O),
    .loops_stencil_valid_ranges_5(loops_stencil_valid_ranges_5_inst0_O),
    .strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr_inst0_O),
    .strg_ub_sram_only_input_addr_gen_0_strides_0(strg_ub_sram_only_input_addr_gen_0_strides_0_inst0_O),
    .strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0(strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0_inst0_O),
    .strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0(strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0_inst0_O),
    .stencil_valid_sched_gen_sched_addr_gen_strides_2(stencil_valid_sched_gen_sched_addr_gen_strides_2_inst0_O),
    .strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr_inst0_O),
    .strg_ub_tb_only_loops_buf2out_read_1_ranges_2(strg_ub_tb_only_loops_buf2out_read_1_ranges_2_inst0_O),
    .loops_stencil_valid_dimensionality(loops_stencil_valid_dimensionality_inst0_O),
    .stencil_valid(LakeTop_W_inst0_stencil_valid),
    .stencil_valid_sched_gen_sched_addr_gen_strides_4(stencil_valid_sched_gen_sched_addr_gen_strides_4_inst0_O),
    .strg_ub_tb_only_tb_read_addr_gen_1_strides_2(strg_ub_tb_only_tb_read_addr_gen_1_strides_2_inst0_O),
    .strg_ub_tb_only_loops_buf2out_read_0_ranges_2(strg_ub_tb_only_loops_buf2out_read_0_ranges_2_inst0_O),
    .strg_ub_tb_only_tb_read_addr_gen_0_strides_0(strg_ub_tb_only_tb_read_addr_gen_0_strides_0_inst0_O),
    .strg_ub_tb_only_loops_buf2out_read_1_ranges_0(strg_ub_tb_only_loops_buf2out_read_1_ranges_0_inst0_O),
    .strg_ub_sram_only_output_addr_gen_1_strides_2(strg_ub_sram_only_output_addr_gen_1_strides_2_inst0_O),
    .strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5(strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5_inst0_O),
    .config_addr_in(OR_config_addr_FEATURE_O),
    .strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr(strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr_inst0_O),
    .strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0(strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0_inst0_O),
    .strg_ub_agg_only_agg_write_addr_gen_0_strides_4(strg_ub_agg_only_agg_write_addr_gen_0_strides_4_inst0_O),
    .strg_ub_tb_only_loops_buf2out_read_0_ranges_1(strg_ub_tb_only_loops_buf2out_read_0_ranges_1_inst0_O),
    .strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5_inst0_O),
    .strg_ub_tb_only_loops_buf2out_read_1_ranges_3(strg_ub_tb_only_loops_buf2out_read_1_ranges_3_inst0_O),
    .strg_ub_agg_only_agg_read_addr_gen_1_strides_5(strg_ub_agg_only_agg_read_addr_gen_1_strides_5_inst0_O),
    .stencil_valid_sched_gen_sched_addr_gen_strides_5(stencil_valid_sched_gen_sched_addr_gen_strides_5_inst0_O),
    .strg_ub_tb_only_tb_write_addr_gen_1_strides_2(strg_ub_tb_only_tb_write_addr_gen_1_strides_2_inst0_O),
    .data_out_0(LakeTop_W_inst0_data_out_0),
    .strg_ub_tb_only_loops_buf2out_read_0_ranges_5(strg_ub_tb_only_loops_buf2out_read_0_ranges_5_inst0_O),
    .strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0(strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0_inst0_O),
    .strg_ub_agg_only_loops_in2buf_1_ranges_0(strg_ub_agg_only_loops_in2buf_1_ranges_0_inst0_O),
    .strg_ub_tb_only_loops_buf2out_read_1_ranges_5(strg_ub_tb_only_loops_buf2out_read_1_ranges_5_inst0_O),
    .strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1(strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1_inst0_O),
    .strg_ub_sram_only_output_addr_gen_0_strides_0(strg_ub_sram_only_output_addr_gen_0_strides_0_inst0_O),
    .strg_ub_tb_only_loops_buf2out_read_0_ranges_0(strg_ub_tb_only_loops_buf2out_read_0_ranges_0_inst0_O),
    .strg_ub_tb_only_tb_read_addr_gen_0_strides_1(strg_ub_tb_only_tb_read_addr_gen_0_strides_1_inst0_O),
    .strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2_inst0_O),
    .strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3(strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3_inst0_O),
    .strg_ub_agg_only_agg_read_addr_gen_1_strides_3(strg_ub_agg_only_agg_read_addr_gen_1_strides_3_inst0_O),
    .strg_ub_tb_only_tb_write_addr_gen_0_strides_1(strg_ub_tb_only_tb_write_addr_gen_0_strides_1_inst0_O),
    .strg_ub_agg_only_loops_in2buf_1_ranges_2(strg_ub_agg_only_loops_in2buf_1_ranges_2_inst0_O),
    .strg_ub_tb_only_tb_write_addr_gen_1_strides_1(strg_ub_tb_only_tb_write_addr_gen_1_strides_1_inst0_O),
    .strg_ub_tb_only_tb_read_addr_gen_1_strides_1(strg_ub_tb_only_tb_read_addr_gen_1_strides_1_inst0_O),
    .stencil_valid_sched_gen_sched_addr_gen_strides_1(stencil_valid_sched_gen_sched_addr_gen_strides_1_inst0_O),
    .strg_ub_sram_only_output_addr_gen_0_strides_1(strg_ub_sram_only_output_addr_gen_0_strides_1_inst0_O),
    .strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr_inst0_O),
    .strg_ub_agg_only_agg_write_addr_gen_0_starting_addr(strg_ub_agg_only_agg_write_addr_gen_0_starting_addr_inst0_O),
    .config_data_in(OR_config_data_FEATURE_O),
    .strg_ub_agg_only_loops_in2buf_1_dimensionality(strg_ub_agg_only_loops_in2buf_1_dimensionality_inst0_O),
    .config_write(OR_CONFIG_RD_SRAM_out),
    .strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5(strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5_inst0_O),
    .strg_ub_agg_only_loops_in2buf_1_ranges_5(strg_ub_agg_only_loops_in2buf_1_ranges_5_inst0_O),
    .strg_ub_agg_only_loops_in2buf_0_ranges_2(strg_ub_agg_only_loops_in2buf_0_ranges_2_inst0_O),
    .strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3(strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3_inst0_O),
    .chain_data_in_1(chain_data_in_1),
    .strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0(strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0_inst0_O),
    .strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2(strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2_inst0_O),
    .strg_ub_tb_only_tb_read_addr_gen_1_strides_5(strg_ub_tb_only_tb_read_addr_gen_1_strides_5_inst0_O),
    .strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0(strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0_inst0_O),
    .strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality_inst0_O),
    .strg_ub_tb_only_tb_read_addr_gen_1_strides_0(strg_ub_tb_only_tb_read_addr_gen_1_strides_0_inst0_O),
    .strg_ub_agg_only_agg_read_addr_gen_1_strides_4(strg_ub_agg_only_agg_read_addr_gen_1_strides_4_inst0_O),
    .strg_ub_agg_only_loops_in2buf_0_dimensionality(strg_ub_agg_only_loops_in2buf_0_dimensionality_inst0_O),
    .strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr_inst0_O),
    .strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5(strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5_inst0_O),
    .strg_ub_agg_only_agg_read_addr_gen_1_starting_addr(strg_ub_agg_only_agg_read_addr_gen_1_starting_addr_inst0_O),
    .config_en(LakeTop_W_inst0_config_en),
    .strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4_inst0_O),
    .strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4_inst0_O),
    .strg_ub_tb_only_tb_read_addr_gen_0_strides_2(strg_ub_tb_only_tb_read_addr_gen_0_strides_2_inst0_O),
    .strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1_inst0_O),
    .strg_ub_tb_only_loops_buf2out_read_0_ranges_4(strg_ub_tb_only_loops_buf2out_read_0_ranges_4_inst0_O),
    .strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2(strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2_inst0_O),
    .strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3_inst0_O),
    .strg_ub_tb_only_tb_write_addr_gen_1_strides_4(strg_ub_tb_only_tb_write_addr_gen_1_strides_4_inst0_O),
    .valid_out(LakeTop_W_inst0_valid_out),
    .strg_ub_tb_only_tb_write_addr_gen_0_strides_5(strg_ub_tb_only_tb_write_addr_gen_0_strides_5_inst0_O),
    .strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality_inst0_O),
    .strg_ub_agg_only_agg_read_addr_gen_0_strides_0(strg_ub_agg_only_agg_read_addr_gen_0_strides_0_inst0_O),
    .strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4(strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4_inst0_O),
    .chain_data_in_0(chain_data_in_0),
    .strg_ub_sram_only_output_addr_gen_0_strides_4(strg_ub_sram_only_output_addr_gen_0_strides_4_inst0_O),
    .strg_ub_agg_only_loops_in2buf_0_ranges_5(strg_ub_agg_only_loops_in2buf_0_ranges_5_inst0_O),
    .strg_ub_tb_only_tb_read_addr_gen_1_strides_3(strg_ub_tb_only_tb_read_addr_gen_1_strides_3_inst0_O),
    .full(LakeTop_W_inst0_full),
    .strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr(strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr_inst0_O),
    .strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3_inst0_O),
    .stencil_valid_sched_gen_sched_addr_gen_strides_3(stencil_valid_sched_gen_sched_addr_gen_strides_3_inst0_O),
    .strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2(strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2_inst0_O),
    .strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5(strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5_inst0_O),
    .strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0_inst0_O),
    .strg_ub_tb_only_loops_buf2out_read_1_ranges_4(strg_ub_tb_only_loops_buf2out_read_1_ranges_4_inst0_O),
    .addr_in_0(addr_in_0),
    .strg_ub_tb_only_tb_read_addr_gen_0_strides_3(strg_ub_tb_only_tb_read_addr_gen_0_strides_3_inst0_O),
    .strg_ub_agg_only_loops_in2buf_1_ranges_4(strg_ub_agg_only_loops_in2buf_1_ranges_4_inst0_O),
    .strg_ub_tb_only_tb_write_addr_gen_0_strides_3(strg_ub_tb_only_tb_write_addr_gen_0_strides_3_inst0_O),
    .strg_ub_tb_only_tb_write_addr_gen_1_strides_5(strg_ub_tb_only_tb_write_addr_gen_1_strides_5_inst0_O),
    .strg_ub_agg_sram_shared_agg_read_sched_gen_0_enable(strg_ub_agg_sram_shared_agg_read_sched_gen_0_enable_inst0_O),
    .strg_ub_agg_only_agg_write_sched_gen_1_enable(strg_ub_agg_only_agg_write_sched_gen_1_enable_inst0_O),
    .fifo_ctrl_fifo_depth(fifo_ctrl_fifo_depth_inst0_O),
    .strg_ub_agg_only_agg_read_addr_gen_0_strides_3(strg_ub_agg_only_agg_read_addr_gen_0_strides_3_inst0_O),
    .strg_ub_tb_only_tb_read_addr_gen_0_strides_4(strg_ub_tb_only_tb_read_addr_gen_0_strides_4_inst0_O),
    .config_read(OR_CONFIG_WR_SRAM_out),
    .strg_ub_tb_only_tb_read_addr_gen_1_strides_4(strg_ub_tb_only_tb_read_addr_gen_1_strides_4_inst0_O),
    .strg_ub_tb_only_tb_write_addr_gen_1_starting_addr(strg_ub_tb_only_tb_write_addr_gen_1_starting_addr_inst0_O),
    .strg_ub_sram_tb_shared_output_sched_gen_0_enable(strg_ub_sram_tb_shared_output_sched_gen_0_enable_inst0_O),
    .strg_ub_tb_only_tb_read_addr_gen_0_starting_addr(strg_ub_tb_only_tb_read_addr_gen_0_starting_addr_inst0_O),
    .strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3(strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3_inst0_O),
    .strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4(strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4_inst0_O),
    .strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0_inst0_O),
    .config_data_out_0(LakeTop_W_inst0_config_data_out_0),
    .strg_ub_agg_only_agg_write_addr_gen_1_strides_5(strg_ub_agg_only_agg_write_addr_gen_1_strides_5_inst0_O),
    .strg_ub_agg_only_agg_write_addr_gen_1_strides_4(strg_ub_agg_only_agg_write_addr_gen_1_strides_4_inst0_O)
);
commonlib_muxn__N84__width32 MuxWrapper_84_32_inst0$Mux84x32_inst0$coreir_commonlib_mux84x32_inst0 (
    .in_data_0(ZextWrapper_23_32_inst0$self_O_in),
    .in_data_1(config_reg_1_O),
    .in_data_10(config_reg_10_O),
    .in_data_11(ZextWrapper_17_32_inst0$self_O_in),
    .in_data_12(config_reg_12_O),
    .in_data_13(config_reg_13_O),
    .in_data_14(config_reg_14_O),
    .in_data_15(ZextWrapper_17_32_inst1$self_O_in),
    .in_data_16(config_reg_16_O),
    .in_data_17(config_reg_17_O),
    .in_data_18(config_reg_18_O),
    .in_data_19(ZextWrapper_20_32_inst0$self_O_in),
    .in_data_2(config_reg_2_O),
    .in_data_20(config_reg_20_O),
    .in_data_21(config_reg_21_O),
    .in_data_22(config_reg_22_O),
    .in_data_23(ZextWrapper_20_32_inst1$self_O_in),
    .in_data_24(config_reg_24_O),
    .in_data_25(config_reg_25_O),
    .in_data_26(ZextWrapper_17_32_inst2$self_O_in),
    .in_data_27(config_reg_27_O),
    .in_data_28(config_reg_28_O),
    .in_data_29(config_reg_29_O),
    .in_data_3(config_reg_3_O),
    .in_data_30(ZextWrapper_17_32_inst3$self_O_in),
    .in_data_31(config_reg_31_O),
    .in_data_32(config_reg_32_O),
    .in_data_33(config_reg_33_O),
    .in_data_34(ZextWrapper_20_32_inst2$self_O_in),
    .in_data_35(config_reg_35_O),
    .in_data_36(config_reg_36_O),
    .in_data_37(config_reg_37_O),
    .in_data_38(ZextWrapper_20_32_inst3$self_O_in),
    .in_data_39(config_reg_39_O),
    .in_data_4(ZextWrapper_23_32_inst1$self_O_in),
    .in_data_40(config_reg_40_O),
    .in_data_41(ZextWrapper_25_32_inst0$self_O_in),
    .in_data_42(ZextWrapper_27_32_inst0$self_O_in),
    .in_data_43(ZextWrapper_27_32_inst1$self_O_in),
    .in_data_44(ZextWrapper_27_32_inst2$self_O_in),
    .in_data_45(ZextWrapper_27_32_inst3$self_O_in),
    .in_data_46(ZextWrapper_27_32_inst4$self_O_in),
    .in_data_47(ZextWrapper_27_32_inst5$self_O_in),
    .in_data_48(ZextWrapper_27_32_inst6$self_O_in),
    .in_data_49(ZextWrapper_27_32_inst7$self_O_in),
    .in_data_5(config_reg_5_O),
    .in_data_50(ZextWrapper_31_32_inst0$self_O_in),
    .in_data_51(config_reg_51_O),
    .in_data_52(config_reg_52_O),
    .in_data_53(config_reg_53_O),
    .in_data_54(ZextWrapper_20_32_inst4$self_O_in),
    .in_data_55(config_reg_55_O),
    .in_data_56(config_reg_56_O),
    .in_data_57(ZextWrapper_17_32_inst4$self_O_in),
    .in_data_58(config_reg_58_O),
    .in_data_59(config_reg_59_O),
    .in_data_6(config_reg_6_O),
    .in_data_60(config_reg_60_O),
    .in_data_61(ZextWrapper_17_32_inst5$self_O_in),
    .in_data_62(config_reg_62_O),
    .in_data_63(config_reg_63_O),
    .in_data_64(config_reg_64_O),
    .in_data_65(ZextWrapper_20_32_inst5$self_O_in),
    .in_data_66(config_reg_66_O),
    .in_data_67(config_reg_67_O),
    .in_data_68(config_reg_68_O),
    .in_data_69(ZextWrapper_20_32_inst6$self_O_in),
    .in_data_7(config_reg_7_O),
    .in_data_70(config_reg_70_O),
    .in_data_71(config_reg_71_O),
    .in_data_72(config_reg_72_O),
    .in_data_73(config_reg_73_O),
    .in_data_74(ZextWrapper_25_32_inst1$self_O_in),
    .in_data_75(config_reg_75_O),
    .in_data_76(config_reg_76_O),
    .in_data_77(config_reg_77_O),
    .in_data_78(ZextWrapper_17_32_inst6$self_O_in),
    .in_data_79(config_reg_79_O),
    .in_data_8(config_reg_8_O),
    .in_data_80(config_reg_80_O),
    .in_data_81(config_reg_81_O),
    .in_data_82(config_reg_82_O),
    .in_data_83(ZextWrapper_29_32_inst0$self_O_in),
    .in_data_9(config_reg_9_O),
    .in_sel(MuxWrapper_84_32_inst0_S_in),
    .out(MuxWrapper_84_32_inst0$Mux84x32_inst0$coreir_commonlib_mux84x32_inst0_out)
);
mantle_wire__typeBitIn7 MuxWrapper_84_32_inst0_S (
    .in(MuxWrapper_84_32_inst0_S_in),
    .out(self_config_config_addr_out[6:0])
);
coreir_or #(
    .width(1)
) OR_CONFIG_EN_SRAM_0 (
    .in0(config_1_write),
    .in1(config_1_read),
    .out(OR_CONFIG_EN_SRAM_0_out)
);
coreir_or #(
    .width(1)
) OR_CONFIG_EN_SRAM_1 (
    .in0(config_2_write),
    .in1(config_2_read),
    .out(OR_CONFIG_EN_SRAM_1_out)
);
coreir_or #(
    .width(1)
) OR_CONFIG_RD_SRAM (
    .in0(config_1_write),
    .in1(config_2_write),
    .out(OR_CONFIG_RD_SRAM_out)
);
coreir_or #(
    .width(1)
) OR_CONFIG_WR_SRAM (
    .in0(config_1_read),
    .in1(config_2_read),
    .out(OR_CONFIG_WR_SRAM_out)
);
Or3x8 OR_config_addr_FEATURE (
    .I0(config_config_addr),
    .I1(config_1_config_addr),
    .I2(config_2_config_addr),
    .O(OR_config_addr_FEATURE_O)
);
Or3x32 OR_config_data_FEATURE (
    .I0(config_config_data),
    .I1(config_1_config_data),
    .I2(config_2_config_data),
    .O(OR_config_data_FEATURE_O)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_17_32_inst0$bit_const_0_None (
    .out(ZextWrapper_17_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit17 ZextWrapper_17_32_inst0$self_I (
    .in(config_reg_11_O),
    .out(ZextWrapper_17_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_17_32_inst0$self_O_out;
assign ZextWrapper_17_32_inst0$self_O_out = {ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$bit_const_0_None_out,ZextWrapper_17_32_inst0$self_I_out[16:0]};
mantle_wire__typeBitIn32 ZextWrapper_17_32_inst0$self_O (
    .in(ZextWrapper_17_32_inst0$self_O_in),
    .out(ZextWrapper_17_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_17_32_inst1$bit_const_0_None (
    .out(ZextWrapper_17_32_inst1$bit_const_0_None_out)
);
mantle_wire__typeBit17 ZextWrapper_17_32_inst1$self_I (
    .in(config_reg_15_O),
    .out(ZextWrapper_17_32_inst1$self_I_out)
);
wire [31:0] ZextWrapper_17_32_inst1$self_O_out;
assign ZextWrapper_17_32_inst1$self_O_out = {ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$bit_const_0_None_out,ZextWrapper_17_32_inst1$self_I_out[16:0]};
mantle_wire__typeBitIn32 ZextWrapper_17_32_inst1$self_O (
    .in(ZextWrapper_17_32_inst1$self_O_in),
    .out(ZextWrapper_17_32_inst1$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_17_32_inst2$bit_const_0_None (
    .out(ZextWrapper_17_32_inst2$bit_const_0_None_out)
);
mantle_wire__typeBit17 ZextWrapper_17_32_inst2$self_I (
    .in(config_reg_26_O),
    .out(ZextWrapper_17_32_inst2$self_I_out)
);
wire [31:0] ZextWrapper_17_32_inst2$self_O_out;
assign ZextWrapper_17_32_inst2$self_O_out = {ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$bit_const_0_None_out,ZextWrapper_17_32_inst2$self_I_out[16:0]};
mantle_wire__typeBitIn32 ZextWrapper_17_32_inst2$self_O (
    .in(ZextWrapper_17_32_inst2$self_O_in),
    .out(ZextWrapper_17_32_inst2$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_17_32_inst3$bit_const_0_None (
    .out(ZextWrapper_17_32_inst3$bit_const_0_None_out)
);
mantle_wire__typeBit17 ZextWrapper_17_32_inst3$self_I (
    .in(config_reg_30_O),
    .out(ZextWrapper_17_32_inst3$self_I_out)
);
wire [31:0] ZextWrapper_17_32_inst3$self_O_out;
assign ZextWrapper_17_32_inst3$self_O_out = {ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$bit_const_0_None_out,ZextWrapper_17_32_inst3$self_I_out[16:0]};
mantle_wire__typeBitIn32 ZextWrapper_17_32_inst3$self_O (
    .in(ZextWrapper_17_32_inst3$self_O_in),
    .out(ZextWrapper_17_32_inst3$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_17_32_inst4$bit_const_0_None (
    .out(ZextWrapper_17_32_inst4$bit_const_0_None_out)
);
mantle_wire__typeBit17 ZextWrapper_17_32_inst4$self_I (
    .in(config_reg_57_O),
    .out(ZextWrapper_17_32_inst4$self_I_out)
);
wire [31:0] ZextWrapper_17_32_inst4$self_O_out;
assign ZextWrapper_17_32_inst4$self_O_out = {ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$bit_const_0_None_out,ZextWrapper_17_32_inst4$self_I_out[16:0]};
mantle_wire__typeBitIn32 ZextWrapper_17_32_inst4$self_O (
    .in(ZextWrapper_17_32_inst4$self_O_in),
    .out(ZextWrapper_17_32_inst4$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_17_32_inst5$bit_const_0_None (
    .out(ZextWrapper_17_32_inst5$bit_const_0_None_out)
);
mantle_wire__typeBit17 ZextWrapper_17_32_inst5$self_I (
    .in(config_reg_61_O),
    .out(ZextWrapper_17_32_inst5$self_I_out)
);
wire [31:0] ZextWrapper_17_32_inst5$self_O_out;
assign ZextWrapper_17_32_inst5$self_O_out = {ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$bit_const_0_None_out,ZextWrapper_17_32_inst5$self_I_out[16:0]};
mantle_wire__typeBitIn32 ZextWrapper_17_32_inst5$self_O (
    .in(ZextWrapper_17_32_inst5$self_O_in),
    .out(ZextWrapper_17_32_inst5$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_17_32_inst6$bit_const_0_None (
    .out(ZextWrapper_17_32_inst6$bit_const_0_None_out)
);
mantle_wire__typeBit17 ZextWrapper_17_32_inst6$self_I (
    .in(config_reg_78_O),
    .out(ZextWrapper_17_32_inst6$self_I_out)
);
wire [31:0] ZextWrapper_17_32_inst6$self_O_out;
assign ZextWrapper_17_32_inst6$self_O_out = {ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$bit_const_0_None_out,ZextWrapper_17_32_inst6$self_I_out[16:0]};
mantle_wire__typeBitIn32 ZextWrapper_17_32_inst6$self_O (
    .in(ZextWrapper_17_32_inst6$self_O_in),
    .out(ZextWrapper_17_32_inst6$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_20_32_inst0$bit_const_0_None (
    .out(ZextWrapper_20_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit20 ZextWrapper_20_32_inst0$self_I (
    .in(config_reg_19_O),
    .out(ZextWrapper_20_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_20_32_inst0$self_O_out;
assign ZextWrapper_20_32_inst0$self_O_out = {ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$bit_const_0_None_out,ZextWrapper_20_32_inst0$self_I_out[19:0]};
mantle_wire__typeBitIn32 ZextWrapper_20_32_inst0$self_O (
    .in(ZextWrapper_20_32_inst0$self_O_in),
    .out(ZextWrapper_20_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_20_32_inst1$bit_const_0_None (
    .out(ZextWrapper_20_32_inst1$bit_const_0_None_out)
);
mantle_wire__typeBit20 ZextWrapper_20_32_inst1$self_I (
    .in(config_reg_23_O),
    .out(ZextWrapper_20_32_inst1$self_I_out)
);
wire [31:0] ZextWrapper_20_32_inst1$self_O_out;
assign ZextWrapper_20_32_inst1$self_O_out = {ZextWrapper_20_32_inst1$bit_const_0_None_out,ZextWrapper_20_32_inst1$bit_const_0_None_out,ZextWrapper_20_32_inst1$bit_const_0_None_out,ZextWrapper_20_32_inst1$bit_const_0_None_out,ZextWrapper_20_32_inst1$bit_const_0_None_out,ZextWrapper_20_32_inst1$bit_const_0_None_out,ZextWrapper_20_32_inst1$bit_const_0_None_out,ZextWrapper_20_32_inst1$bit_const_0_None_out,ZextWrapper_20_32_inst1$bit_const_0_None_out,ZextWrapper_20_32_inst1$bit_const_0_None_out,ZextWrapper_20_32_inst1$bit_const_0_None_out,ZextWrapper_20_32_inst1$bit_const_0_None_out,ZextWrapper_20_32_inst1$self_I_out[19:0]};
mantle_wire__typeBitIn32 ZextWrapper_20_32_inst1$self_O (
    .in(ZextWrapper_20_32_inst1$self_O_in),
    .out(ZextWrapper_20_32_inst1$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_20_32_inst2$bit_const_0_None (
    .out(ZextWrapper_20_32_inst2$bit_const_0_None_out)
);
mantle_wire__typeBit20 ZextWrapper_20_32_inst2$self_I (
    .in(config_reg_34_O),
    .out(ZextWrapper_20_32_inst2$self_I_out)
);
wire [31:0] ZextWrapper_20_32_inst2$self_O_out;
assign ZextWrapper_20_32_inst2$self_O_out = {ZextWrapper_20_32_inst2$bit_const_0_None_out,ZextWrapper_20_32_inst2$bit_const_0_None_out,ZextWrapper_20_32_inst2$bit_const_0_None_out,ZextWrapper_20_32_inst2$bit_const_0_None_out,ZextWrapper_20_32_inst2$bit_const_0_None_out,ZextWrapper_20_32_inst2$bit_const_0_None_out,ZextWrapper_20_32_inst2$bit_const_0_None_out,ZextWrapper_20_32_inst2$bit_const_0_None_out,ZextWrapper_20_32_inst2$bit_const_0_None_out,ZextWrapper_20_32_inst2$bit_const_0_None_out,ZextWrapper_20_32_inst2$bit_const_0_None_out,ZextWrapper_20_32_inst2$bit_const_0_None_out,ZextWrapper_20_32_inst2$self_I_out[19:0]};
mantle_wire__typeBitIn32 ZextWrapper_20_32_inst2$self_O (
    .in(ZextWrapper_20_32_inst2$self_O_in),
    .out(ZextWrapper_20_32_inst2$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_20_32_inst3$bit_const_0_None (
    .out(ZextWrapper_20_32_inst3$bit_const_0_None_out)
);
mantle_wire__typeBit20 ZextWrapper_20_32_inst3$self_I (
    .in(config_reg_38_O),
    .out(ZextWrapper_20_32_inst3$self_I_out)
);
wire [31:0] ZextWrapper_20_32_inst3$self_O_out;
assign ZextWrapper_20_32_inst3$self_O_out = {ZextWrapper_20_32_inst3$bit_const_0_None_out,ZextWrapper_20_32_inst3$bit_const_0_None_out,ZextWrapper_20_32_inst3$bit_const_0_None_out,ZextWrapper_20_32_inst3$bit_const_0_None_out,ZextWrapper_20_32_inst3$bit_const_0_None_out,ZextWrapper_20_32_inst3$bit_const_0_None_out,ZextWrapper_20_32_inst3$bit_const_0_None_out,ZextWrapper_20_32_inst3$bit_const_0_None_out,ZextWrapper_20_32_inst3$bit_const_0_None_out,ZextWrapper_20_32_inst3$bit_const_0_None_out,ZextWrapper_20_32_inst3$bit_const_0_None_out,ZextWrapper_20_32_inst3$bit_const_0_None_out,ZextWrapper_20_32_inst3$self_I_out[19:0]};
mantle_wire__typeBitIn32 ZextWrapper_20_32_inst3$self_O (
    .in(ZextWrapper_20_32_inst3$self_O_in),
    .out(ZextWrapper_20_32_inst3$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_20_32_inst4$bit_const_0_None (
    .out(ZextWrapper_20_32_inst4$bit_const_0_None_out)
);
mantle_wire__typeBit20 ZextWrapper_20_32_inst4$self_I (
    .in(config_reg_54_O),
    .out(ZextWrapper_20_32_inst4$self_I_out)
);
wire [31:0] ZextWrapper_20_32_inst4$self_O_out;
assign ZextWrapper_20_32_inst4$self_O_out = {ZextWrapper_20_32_inst4$bit_const_0_None_out,ZextWrapper_20_32_inst4$bit_const_0_None_out,ZextWrapper_20_32_inst4$bit_const_0_None_out,ZextWrapper_20_32_inst4$bit_const_0_None_out,ZextWrapper_20_32_inst4$bit_const_0_None_out,ZextWrapper_20_32_inst4$bit_const_0_None_out,ZextWrapper_20_32_inst4$bit_const_0_None_out,ZextWrapper_20_32_inst4$bit_const_0_None_out,ZextWrapper_20_32_inst4$bit_const_0_None_out,ZextWrapper_20_32_inst4$bit_const_0_None_out,ZextWrapper_20_32_inst4$bit_const_0_None_out,ZextWrapper_20_32_inst4$bit_const_0_None_out,ZextWrapper_20_32_inst4$self_I_out[19:0]};
mantle_wire__typeBitIn32 ZextWrapper_20_32_inst4$self_O (
    .in(ZextWrapper_20_32_inst4$self_O_in),
    .out(ZextWrapper_20_32_inst4$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_20_32_inst5$bit_const_0_None (
    .out(ZextWrapper_20_32_inst5$bit_const_0_None_out)
);
mantle_wire__typeBit20 ZextWrapper_20_32_inst5$self_I (
    .in(config_reg_65_O),
    .out(ZextWrapper_20_32_inst5$self_I_out)
);
wire [31:0] ZextWrapper_20_32_inst5$self_O_out;
assign ZextWrapper_20_32_inst5$self_O_out = {ZextWrapper_20_32_inst5$bit_const_0_None_out,ZextWrapper_20_32_inst5$bit_const_0_None_out,ZextWrapper_20_32_inst5$bit_const_0_None_out,ZextWrapper_20_32_inst5$bit_const_0_None_out,ZextWrapper_20_32_inst5$bit_const_0_None_out,ZextWrapper_20_32_inst5$bit_const_0_None_out,ZextWrapper_20_32_inst5$bit_const_0_None_out,ZextWrapper_20_32_inst5$bit_const_0_None_out,ZextWrapper_20_32_inst5$bit_const_0_None_out,ZextWrapper_20_32_inst5$bit_const_0_None_out,ZextWrapper_20_32_inst5$bit_const_0_None_out,ZextWrapper_20_32_inst5$bit_const_0_None_out,ZextWrapper_20_32_inst5$self_I_out[19:0]};
mantle_wire__typeBitIn32 ZextWrapper_20_32_inst5$self_O (
    .in(ZextWrapper_20_32_inst5$self_O_in),
    .out(ZextWrapper_20_32_inst5$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_20_32_inst6$bit_const_0_None (
    .out(ZextWrapper_20_32_inst6$bit_const_0_None_out)
);
mantle_wire__typeBit20 ZextWrapper_20_32_inst6$self_I (
    .in(config_reg_69_O),
    .out(ZextWrapper_20_32_inst6$self_I_out)
);
wire [31:0] ZextWrapper_20_32_inst6$self_O_out;
assign ZextWrapper_20_32_inst6$self_O_out = {ZextWrapper_20_32_inst6$bit_const_0_None_out,ZextWrapper_20_32_inst6$bit_const_0_None_out,ZextWrapper_20_32_inst6$bit_const_0_None_out,ZextWrapper_20_32_inst6$bit_const_0_None_out,ZextWrapper_20_32_inst6$bit_const_0_None_out,ZextWrapper_20_32_inst6$bit_const_0_None_out,ZextWrapper_20_32_inst6$bit_const_0_None_out,ZextWrapper_20_32_inst6$bit_const_0_None_out,ZextWrapper_20_32_inst6$bit_const_0_None_out,ZextWrapper_20_32_inst6$bit_const_0_None_out,ZextWrapper_20_32_inst6$bit_const_0_None_out,ZextWrapper_20_32_inst6$bit_const_0_None_out,ZextWrapper_20_32_inst6$self_I_out[19:0]};
mantle_wire__typeBitIn32 ZextWrapper_20_32_inst6$self_O (
    .in(ZextWrapper_20_32_inst6$self_O_in),
    .out(ZextWrapper_20_32_inst6$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_23_32_inst0$bit_const_0_None (
    .out(ZextWrapper_23_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit23 ZextWrapper_23_32_inst0$self_I (
    .in(config_reg_0_O),
    .out(ZextWrapper_23_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_23_32_inst0$self_O_out;
assign ZextWrapper_23_32_inst0$self_O_out = {ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$bit_const_0_None_out,ZextWrapper_23_32_inst0$self_I_out[22:0]};
mantle_wire__typeBitIn32 ZextWrapper_23_32_inst0$self_O (
    .in(ZextWrapper_23_32_inst0$self_O_in),
    .out(ZextWrapper_23_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_23_32_inst1$bit_const_0_None (
    .out(ZextWrapper_23_32_inst1$bit_const_0_None_out)
);
mantle_wire__typeBit23 ZextWrapper_23_32_inst1$self_I (
    .in(config_reg_4_O),
    .out(ZextWrapper_23_32_inst1$self_I_out)
);
wire [31:0] ZextWrapper_23_32_inst1$self_O_out;
assign ZextWrapper_23_32_inst1$self_O_out = {ZextWrapper_23_32_inst1$bit_const_0_None_out,ZextWrapper_23_32_inst1$bit_const_0_None_out,ZextWrapper_23_32_inst1$bit_const_0_None_out,ZextWrapper_23_32_inst1$bit_const_0_None_out,ZextWrapper_23_32_inst1$bit_const_0_None_out,ZextWrapper_23_32_inst1$bit_const_0_None_out,ZextWrapper_23_32_inst1$bit_const_0_None_out,ZextWrapper_23_32_inst1$bit_const_0_None_out,ZextWrapper_23_32_inst1$bit_const_0_None_out,ZextWrapper_23_32_inst1$self_I_out[22:0]};
mantle_wire__typeBitIn32 ZextWrapper_23_32_inst1$self_O (
    .in(ZextWrapper_23_32_inst1$self_O_in),
    .out(ZextWrapper_23_32_inst1$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_25_32_inst0$bit_const_0_None (
    .out(ZextWrapper_25_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit25 ZextWrapper_25_32_inst0$self_I (
    .in(config_reg_41_O),
    .out(ZextWrapper_25_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_25_32_inst0$self_O_out;
assign ZextWrapper_25_32_inst0$self_O_out = {ZextWrapper_25_32_inst0$bit_const_0_None_out,ZextWrapper_25_32_inst0$bit_const_0_None_out,ZextWrapper_25_32_inst0$bit_const_0_None_out,ZextWrapper_25_32_inst0$bit_const_0_None_out,ZextWrapper_25_32_inst0$bit_const_0_None_out,ZextWrapper_25_32_inst0$bit_const_0_None_out,ZextWrapper_25_32_inst0$bit_const_0_None_out,ZextWrapper_25_32_inst0$self_I_out[24:0]};
mantle_wire__typeBitIn32 ZextWrapper_25_32_inst0$self_O (
    .in(ZextWrapper_25_32_inst0$self_O_in),
    .out(ZextWrapper_25_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_25_32_inst1$bit_const_0_None (
    .out(ZextWrapper_25_32_inst1$bit_const_0_None_out)
);
mantle_wire__typeBit25 ZextWrapper_25_32_inst1$self_I (
    .in(config_reg_74_O),
    .out(ZextWrapper_25_32_inst1$self_I_out)
);
wire [31:0] ZextWrapper_25_32_inst1$self_O_out;
assign ZextWrapper_25_32_inst1$self_O_out = {ZextWrapper_25_32_inst1$bit_const_0_None_out,ZextWrapper_25_32_inst1$bit_const_0_None_out,ZextWrapper_25_32_inst1$bit_const_0_None_out,ZextWrapper_25_32_inst1$bit_const_0_None_out,ZextWrapper_25_32_inst1$bit_const_0_None_out,ZextWrapper_25_32_inst1$bit_const_0_None_out,ZextWrapper_25_32_inst1$bit_const_0_None_out,ZextWrapper_25_32_inst1$self_I_out[24:0]};
mantle_wire__typeBitIn32 ZextWrapper_25_32_inst1$self_O (
    .in(ZextWrapper_25_32_inst1$self_O_in),
    .out(ZextWrapper_25_32_inst1$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_27_32_inst0$bit_const_0_None (
    .out(ZextWrapper_27_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit27 ZextWrapper_27_32_inst0$self_I (
    .in(config_reg_42_O),
    .out(ZextWrapper_27_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_27_32_inst0$self_O_out;
assign ZextWrapper_27_32_inst0$self_O_out = {ZextWrapper_27_32_inst0$bit_const_0_None_out,ZextWrapper_27_32_inst0$bit_const_0_None_out,ZextWrapper_27_32_inst0$bit_const_0_None_out,ZextWrapper_27_32_inst0$bit_const_0_None_out,ZextWrapper_27_32_inst0$bit_const_0_None_out,ZextWrapper_27_32_inst0$self_I_out[26:0]};
mantle_wire__typeBitIn32 ZextWrapper_27_32_inst0$self_O (
    .in(ZextWrapper_27_32_inst0$self_O_in),
    .out(ZextWrapper_27_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_27_32_inst1$bit_const_0_None (
    .out(ZextWrapper_27_32_inst1$bit_const_0_None_out)
);
mantle_wire__typeBit27 ZextWrapper_27_32_inst1$self_I (
    .in(config_reg_43_O),
    .out(ZextWrapper_27_32_inst1$self_I_out)
);
wire [31:0] ZextWrapper_27_32_inst1$self_O_out;
assign ZextWrapper_27_32_inst1$self_O_out = {ZextWrapper_27_32_inst1$bit_const_0_None_out,ZextWrapper_27_32_inst1$bit_const_0_None_out,ZextWrapper_27_32_inst1$bit_const_0_None_out,ZextWrapper_27_32_inst1$bit_const_0_None_out,ZextWrapper_27_32_inst1$bit_const_0_None_out,ZextWrapper_27_32_inst1$self_I_out[26:0]};
mantle_wire__typeBitIn32 ZextWrapper_27_32_inst1$self_O (
    .in(ZextWrapper_27_32_inst1$self_O_in),
    .out(ZextWrapper_27_32_inst1$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_27_32_inst2$bit_const_0_None (
    .out(ZextWrapper_27_32_inst2$bit_const_0_None_out)
);
mantle_wire__typeBit27 ZextWrapper_27_32_inst2$self_I (
    .in(config_reg_44_O),
    .out(ZextWrapper_27_32_inst2$self_I_out)
);
wire [31:0] ZextWrapper_27_32_inst2$self_O_out;
assign ZextWrapper_27_32_inst2$self_O_out = {ZextWrapper_27_32_inst2$bit_const_0_None_out,ZextWrapper_27_32_inst2$bit_const_0_None_out,ZextWrapper_27_32_inst2$bit_const_0_None_out,ZextWrapper_27_32_inst2$bit_const_0_None_out,ZextWrapper_27_32_inst2$bit_const_0_None_out,ZextWrapper_27_32_inst2$self_I_out[26:0]};
mantle_wire__typeBitIn32 ZextWrapper_27_32_inst2$self_O (
    .in(ZextWrapper_27_32_inst2$self_O_in),
    .out(ZextWrapper_27_32_inst2$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_27_32_inst3$bit_const_0_None (
    .out(ZextWrapper_27_32_inst3$bit_const_0_None_out)
);
mantle_wire__typeBit27 ZextWrapper_27_32_inst3$self_I (
    .in(config_reg_45_O),
    .out(ZextWrapper_27_32_inst3$self_I_out)
);
wire [31:0] ZextWrapper_27_32_inst3$self_O_out;
assign ZextWrapper_27_32_inst3$self_O_out = {ZextWrapper_27_32_inst3$bit_const_0_None_out,ZextWrapper_27_32_inst3$bit_const_0_None_out,ZextWrapper_27_32_inst3$bit_const_0_None_out,ZextWrapper_27_32_inst3$bit_const_0_None_out,ZextWrapper_27_32_inst3$bit_const_0_None_out,ZextWrapper_27_32_inst3$self_I_out[26:0]};
mantle_wire__typeBitIn32 ZextWrapper_27_32_inst3$self_O (
    .in(ZextWrapper_27_32_inst3$self_O_in),
    .out(ZextWrapper_27_32_inst3$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_27_32_inst4$bit_const_0_None (
    .out(ZextWrapper_27_32_inst4$bit_const_0_None_out)
);
mantle_wire__typeBit27 ZextWrapper_27_32_inst4$self_I (
    .in(config_reg_46_O),
    .out(ZextWrapper_27_32_inst4$self_I_out)
);
wire [31:0] ZextWrapper_27_32_inst4$self_O_out;
assign ZextWrapper_27_32_inst4$self_O_out = {ZextWrapper_27_32_inst4$bit_const_0_None_out,ZextWrapper_27_32_inst4$bit_const_0_None_out,ZextWrapper_27_32_inst4$bit_const_0_None_out,ZextWrapper_27_32_inst4$bit_const_0_None_out,ZextWrapper_27_32_inst4$bit_const_0_None_out,ZextWrapper_27_32_inst4$self_I_out[26:0]};
mantle_wire__typeBitIn32 ZextWrapper_27_32_inst4$self_O (
    .in(ZextWrapper_27_32_inst4$self_O_in),
    .out(ZextWrapper_27_32_inst4$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_27_32_inst5$bit_const_0_None (
    .out(ZextWrapper_27_32_inst5$bit_const_0_None_out)
);
mantle_wire__typeBit27 ZextWrapper_27_32_inst5$self_I (
    .in(config_reg_47_O),
    .out(ZextWrapper_27_32_inst5$self_I_out)
);
wire [31:0] ZextWrapper_27_32_inst5$self_O_out;
assign ZextWrapper_27_32_inst5$self_O_out = {ZextWrapper_27_32_inst5$bit_const_0_None_out,ZextWrapper_27_32_inst5$bit_const_0_None_out,ZextWrapper_27_32_inst5$bit_const_0_None_out,ZextWrapper_27_32_inst5$bit_const_0_None_out,ZextWrapper_27_32_inst5$bit_const_0_None_out,ZextWrapper_27_32_inst5$self_I_out[26:0]};
mantle_wire__typeBitIn32 ZextWrapper_27_32_inst5$self_O (
    .in(ZextWrapper_27_32_inst5$self_O_in),
    .out(ZextWrapper_27_32_inst5$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_27_32_inst6$bit_const_0_None (
    .out(ZextWrapper_27_32_inst6$bit_const_0_None_out)
);
mantle_wire__typeBit27 ZextWrapper_27_32_inst6$self_I (
    .in(config_reg_48_O),
    .out(ZextWrapper_27_32_inst6$self_I_out)
);
wire [31:0] ZextWrapper_27_32_inst6$self_O_out;
assign ZextWrapper_27_32_inst6$self_O_out = {ZextWrapper_27_32_inst6$bit_const_0_None_out,ZextWrapper_27_32_inst6$bit_const_0_None_out,ZextWrapper_27_32_inst6$bit_const_0_None_out,ZextWrapper_27_32_inst6$bit_const_0_None_out,ZextWrapper_27_32_inst6$bit_const_0_None_out,ZextWrapper_27_32_inst6$self_I_out[26:0]};
mantle_wire__typeBitIn32 ZextWrapper_27_32_inst6$self_O (
    .in(ZextWrapper_27_32_inst6$self_O_in),
    .out(ZextWrapper_27_32_inst6$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_27_32_inst7$bit_const_0_None (
    .out(ZextWrapper_27_32_inst7$bit_const_0_None_out)
);
mantle_wire__typeBit27 ZextWrapper_27_32_inst7$self_I (
    .in(config_reg_49_O),
    .out(ZextWrapper_27_32_inst7$self_I_out)
);
wire [31:0] ZextWrapper_27_32_inst7$self_O_out;
assign ZextWrapper_27_32_inst7$self_O_out = {ZextWrapper_27_32_inst7$bit_const_0_None_out,ZextWrapper_27_32_inst7$bit_const_0_None_out,ZextWrapper_27_32_inst7$bit_const_0_None_out,ZextWrapper_27_32_inst7$bit_const_0_None_out,ZextWrapper_27_32_inst7$bit_const_0_None_out,ZextWrapper_27_32_inst7$self_I_out[26:0]};
mantle_wire__typeBitIn32 ZextWrapper_27_32_inst7$self_O (
    .in(ZextWrapper_27_32_inst7$self_O_in),
    .out(ZextWrapper_27_32_inst7$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_29_32_inst0$bit_const_0_None (
    .out(ZextWrapper_29_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit29 ZextWrapper_29_32_inst0$self_I (
    .in(config_reg_83_O),
    .out(ZextWrapper_29_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_29_32_inst0$self_O_out;
assign ZextWrapper_29_32_inst0$self_O_out = {ZextWrapper_29_32_inst0$bit_const_0_None_out,ZextWrapper_29_32_inst0$bit_const_0_None_out,ZextWrapper_29_32_inst0$bit_const_0_None_out,ZextWrapper_29_32_inst0$self_I_out[28:0]};
mantle_wire__typeBitIn32 ZextWrapper_29_32_inst0$self_O (
    .in(ZextWrapper_29_32_inst0$self_O_in),
    .out(ZextWrapper_29_32_inst0$self_O_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_31_32_inst0$bit_const_0_None (
    .out(ZextWrapper_31_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit31 ZextWrapper_31_32_inst0$self_I (
    .in(config_reg_50_O),
    .out(ZextWrapper_31_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_31_32_inst0$self_O_out;
assign ZextWrapper_31_32_inst0$self_O_out = {ZextWrapper_31_32_inst0$bit_const_0_None_out,ZextWrapper_31_32_inst0$self_I_out[30:0]};
mantle_wire__typeBitIn32 ZextWrapper_31_32_inst0$self_O (
    .in(ZextWrapper_31_32_inst0$self_O_in),
    .out(ZextWrapper_31_32_inst0$self_O_out)
);
chain_chain_en chain_chain_en_inst0 (
    .I(config_reg_0_O),
    .O(chain_chain_en_inst0_O)
);
ConfigRegister_23_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_1 config_reg_1 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_1_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_10 config_reg_10 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_10_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_17_8_32_11 config_reg_11 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_11_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_12 config_reg_12 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_12_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_13 config_reg_13 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_13_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_14 config_reg_14 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_14_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_17_8_32_15 config_reg_15 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_15_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_16 config_reg_16 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_16_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_17 config_reg_17 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_17_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_18 config_reg_18 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_18_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_20_8_32_19 config_reg_19 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_19_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_2 config_reg_2 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_2_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_20 config_reg_20 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_20_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_21 config_reg_21 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_21_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_22 config_reg_22 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_22_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_20_8_32_23 config_reg_23 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_23_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_24 config_reg_24 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_24_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_25 config_reg_25 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_25_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_17_8_32_26 config_reg_26 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_26_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_27 config_reg_27 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_27_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_28 config_reg_28 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_28_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_29 config_reg_29 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_29_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_3 config_reg_3 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_3_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_17_8_32_30 config_reg_30 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_30_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_31 config_reg_31 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_31_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_32 config_reg_32 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_32_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_33 config_reg_33 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_33_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_20_8_32_34 config_reg_34 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_34_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_35 config_reg_35 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_35_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_36 config_reg_36 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_36_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_37 config_reg_37 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_37_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_20_8_32_38 config_reg_38 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_38_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_39 config_reg_39 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_39_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_23_8_32_4 config_reg_4 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_4_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_40 config_reg_40 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_40_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_25_8_32_41 config_reg_41 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_41_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_27_8_32_42 config_reg_42 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_42_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_27_8_32_43 config_reg_43 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_43_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_27_8_32_44 config_reg_44 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_44_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_27_8_32_45 config_reg_45 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_45_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_27_8_32_46 config_reg_46 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_46_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_27_8_32_47 config_reg_47 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_47_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_27_8_32_48 config_reg_48 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_48_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_27_8_32_49 config_reg_49 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_49_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_5 config_reg_5 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_5_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_31_8_32_50 config_reg_50 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_50_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_51 config_reg_51 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_51_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_52 config_reg_52 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_52_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_53 config_reg_53 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_53_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_20_8_32_54 config_reg_54 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_54_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_55 config_reg_55 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_55_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_56 config_reg_56 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_56_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_17_8_32_57 config_reg_57 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_57_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_58 config_reg_58 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_58_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_59 config_reg_59 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_59_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_6 config_reg_6 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_6_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_60 config_reg_60 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_60_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_17_8_32_61 config_reg_61 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_61_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_62 config_reg_62 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_62_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_63 config_reg_63 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_63_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_64 config_reg_64 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_64_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_20_8_32_65 config_reg_65 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_65_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_66 config_reg_66 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_66_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_67 config_reg_67 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_67_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_68 config_reg_68 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_68_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_20_8_32_69 config_reg_69 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_69_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_7 config_reg_7 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_7_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_70 config_reg_70 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_70_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_71 config_reg_71 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_71_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_72 config_reg_72 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_72_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_73 config_reg_73 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_73_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_25_8_32_74 config_reg_74 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_74_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_75 config_reg_75 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_75_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_76 config_reg_76 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_76_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_77 config_reg_77 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_77_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_17_8_32_78 config_reg_78 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_78_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_79 config_reg_79 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_79_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_8 config_reg_8 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_8_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_80 config_reg_80 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_80_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_81 config_reg_81 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_81_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_82 config_reg_82 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_82_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_29_8_32_83 config_reg_83 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_83_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_9 config_reg_9 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_9_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
coreir_wrap coreir_wrapInAsyncReset_inst0 (
    .in(reset),
    .out(coreir_wrapInAsyncReset_inst0_out)
);
coreir_wrap coreir_wrapOutAsyncReset_inst0 (
    .in(Invert1_inst0_out[0]),
    .out(coreir_wrapOutAsyncReset_inst0_out)
);
fifo_ctrl_fifo_depth fifo_ctrl_fifo_depth_inst0 (
    .I(config_reg_0_O),
    .O(fifo_ctrl_fifo_depth_inst0_O)
);
flush_reg_sel flush_reg_sel_inst0 (
    .I(config_reg_0_O),
    .O(flush_reg_sel_inst0_O)
);
flush_reg_value flush_reg_value_inst0 (
    .I(config_reg_0_O),
    .O(flush_reg_value_inst0_O)
);
coreir_mux #(
    .width(1)
) flush_sel$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(flush),
    .in1(flush_reg_value_inst0_O),
    .sel(flush_reg_sel_inst0_O[0]),
    .out(flush_sel$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
loops_stencil_valid_dimensionality loops_stencil_valid_dimensionality_inst0 (
    .I(config_reg_0_O),
    .O(loops_stencil_valid_dimensionality_inst0_O)
);
loops_stencil_valid_ranges_0 loops_stencil_valid_ranges_0_inst0 (
    .I(config_reg_1_O),
    .O(loops_stencil_valid_ranges_0_inst0_O)
);
loops_stencil_valid_ranges_1 loops_stencil_valid_ranges_1_inst0 (
    .I(config_reg_1_O),
    .O(loops_stencil_valid_ranges_1_inst0_O)
);
loops_stencil_valid_ranges_2 loops_stencil_valid_ranges_2_inst0 (
    .I(config_reg_2_O),
    .O(loops_stencil_valid_ranges_2_inst0_O)
);
loops_stencil_valid_ranges_3 loops_stencil_valid_ranges_3_inst0 (
    .I(config_reg_2_O),
    .O(loops_stencil_valid_ranges_3_inst0_O)
);
loops_stencil_valid_ranges_4 loops_stencil_valid_ranges_4_inst0 (
    .I(config_reg_3_O),
    .O(loops_stencil_valid_ranges_4_inst0_O)
);
loops_stencil_valid_ranges_5 loops_stencil_valid_ranges_5_inst0 (
    .I(config_reg_3_O),
    .O(loops_stencil_valid_ranges_5_inst0_O)
);
mode mode_inst0 (
    .I(config_reg_4_O),
    .O(mode_inst0_O)
);
ren_in_0_reg_sel ren_in_0_reg_sel_inst0 (
    .I(config_reg_4_O),
    .O(ren_in_0_reg_sel_inst0_O)
);
ren_in_0_reg_value ren_in_0_reg_value_inst0 (
    .I(config_reg_4_O),
    .O(ren_in_0_reg_value_inst0_O)
);
coreir_mux #(
    .width(1)
) ren_in_0_sel$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(ren_in_0),
    .in1(ren_in_0_reg_value_inst0_O),
    .sel(ren_in_0_reg_sel_inst0_O[0]),
    .out(ren_in_0_sel$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
ren_in_1_reg_sel ren_in_1_reg_sel_inst0 (
    .I(config_reg_4_O),
    .O(ren_in_1_reg_sel_inst0_O)
);
ren_in_1_reg_value ren_in_1_reg_value_inst0 (
    .I(config_reg_4_O),
    .O(ren_in_1_reg_value_inst0_O)
);
coreir_mux #(
    .width(1)
) ren_in_1_sel$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(ren_in_1),
    .in1(ren_in_1_reg_value_inst0_O),
    .sel(ren_in_1_reg_sel_inst0_O[0]),
    .out(ren_in_1_sel$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
mantle_wire__typeBit8 self_config_config_addr (
    .in(config_config_addr),
    .out(self_config_config_addr_out)
);
stencil_valid_sched_gen_enable stencil_valid_sched_gen_enable_inst0 (
    .I(config_reg_4_O),
    .O(stencil_valid_sched_gen_enable_inst0_O)
);
stencil_valid_sched_gen_sched_addr_gen_starting_addr stencil_valid_sched_gen_sched_addr_gen_starting_addr_inst0 (
    .I(config_reg_4_O),
    .O(stencil_valid_sched_gen_sched_addr_gen_starting_addr_inst0_O)
);
stencil_valid_sched_gen_sched_addr_gen_strides_0 stencil_valid_sched_gen_sched_addr_gen_strides_0_inst0 (
    .I(config_reg_5_O),
    .O(stencil_valid_sched_gen_sched_addr_gen_strides_0_inst0_O)
);
stencil_valid_sched_gen_sched_addr_gen_strides_1 stencil_valid_sched_gen_sched_addr_gen_strides_1_inst0 (
    .I(config_reg_5_O),
    .O(stencil_valid_sched_gen_sched_addr_gen_strides_1_inst0_O)
);
stencil_valid_sched_gen_sched_addr_gen_strides_2 stencil_valid_sched_gen_sched_addr_gen_strides_2_inst0 (
    .I(config_reg_6_O),
    .O(stencil_valid_sched_gen_sched_addr_gen_strides_2_inst0_O)
);
stencil_valid_sched_gen_sched_addr_gen_strides_3 stencil_valid_sched_gen_sched_addr_gen_strides_3_inst0 (
    .I(config_reg_6_O),
    .O(stencil_valid_sched_gen_sched_addr_gen_strides_3_inst0_O)
);
stencil_valid_sched_gen_sched_addr_gen_strides_4 stencil_valid_sched_gen_sched_addr_gen_strides_4_inst0 (
    .I(config_reg_7_O),
    .O(stencil_valid_sched_gen_sched_addr_gen_strides_4_inst0_O)
);
stencil_valid_sched_gen_sched_addr_gen_strides_5 stencil_valid_sched_gen_sched_addr_gen_strides_5_inst0 (
    .I(config_reg_7_O),
    .O(stencil_valid_sched_gen_sched_addr_gen_strides_5_inst0_O)
);
strg_ub_agg_only_agg_read_addr_gen_0_starting_addr strg_ub_agg_only_agg_read_addr_gen_0_starting_addr_inst0 (
    .I(config_reg_8_O),
    .O(strg_ub_agg_only_agg_read_addr_gen_0_starting_addr_inst0_O)
);
strg_ub_agg_only_agg_read_addr_gen_0_strides_0 strg_ub_agg_only_agg_read_addr_gen_0_strides_0_inst0 (
    .I(config_reg_8_O),
    .O(strg_ub_agg_only_agg_read_addr_gen_0_strides_0_inst0_O)
);
strg_ub_agg_only_agg_read_addr_gen_0_strides_1 strg_ub_agg_only_agg_read_addr_gen_0_strides_1_inst0 (
    .I(config_reg_8_O),
    .O(strg_ub_agg_only_agg_read_addr_gen_0_strides_1_inst0_O)
);
strg_ub_agg_only_agg_read_addr_gen_0_strides_2 strg_ub_agg_only_agg_read_addr_gen_0_strides_2_inst0 (
    .I(config_reg_8_O),
    .O(strg_ub_agg_only_agg_read_addr_gen_0_strides_2_inst0_O)
);
strg_ub_agg_only_agg_read_addr_gen_0_strides_3 strg_ub_agg_only_agg_read_addr_gen_0_strides_3_inst0 (
    .I(config_reg_8_O),
    .O(strg_ub_agg_only_agg_read_addr_gen_0_strides_3_inst0_O)
);
strg_ub_agg_only_agg_read_addr_gen_0_strides_4 strg_ub_agg_only_agg_read_addr_gen_0_strides_4_inst0 (
    .I(config_reg_8_O),
    .O(strg_ub_agg_only_agg_read_addr_gen_0_strides_4_inst0_O)
);
strg_ub_agg_only_agg_read_addr_gen_0_strides_5 strg_ub_agg_only_agg_read_addr_gen_0_strides_5_inst0 (
    .I(config_reg_8_O),
    .O(strg_ub_agg_only_agg_read_addr_gen_0_strides_5_inst0_O)
);
strg_ub_agg_only_agg_read_addr_gen_1_starting_addr strg_ub_agg_only_agg_read_addr_gen_1_starting_addr_inst0 (
    .I(config_reg_8_O),
    .O(strg_ub_agg_only_agg_read_addr_gen_1_starting_addr_inst0_O)
);
strg_ub_agg_only_agg_read_addr_gen_1_strides_0 strg_ub_agg_only_agg_read_addr_gen_1_strides_0_inst0 (
    .I(config_reg_9_O),
    .O(strg_ub_agg_only_agg_read_addr_gen_1_strides_0_inst0_O)
);
strg_ub_agg_only_agg_read_addr_gen_1_strides_1 strg_ub_agg_only_agg_read_addr_gen_1_strides_1_inst0 (
    .I(config_reg_9_O),
    .O(strg_ub_agg_only_agg_read_addr_gen_1_strides_1_inst0_O)
);
strg_ub_agg_only_agg_read_addr_gen_1_strides_2 strg_ub_agg_only_agg_read_addr_gen_1_strides_2_inst0 (
    .I(config_reg_9_O),
    .O(strg_ub_agg_only_agg_read_addr_gen_1_strides_2_inst0_O)
);
strg_ub_agg_only_agg_read_addr_gen_1_strides_3 strg_ub_agg_only_agg_read_addr_gen_1_strides_3_inst0 (
    .I(config_reg_9_O),
    .O(strg_ub_agg_only_agg_read_addr_gen_1_strides_3_inst0_O)
);
strg_ub_agg_only_agg_read_addr_gen_1_strides_4 strg_ub_agg_only_agg_read_addr_gen_1_strides_4_inst0 (
    .I(config_reg_9_O),
    .O(strg_ub_agg_only_agg_read_addr_gen_1_strides_4_inst0_O)
);
strg_ub_agg_only_agg_read_addr_gen_1_strides_5 strg_ub_agg_only_agg_read_addr_gen_1_strides_5_inst0 (
    .I(config_reg_9_O),
    .O(strg_ub_agg_only_agg_read_addr_gen_1_strides_5_inst0_O)
);
strg_ub_agg_only_agg_write_addr_gen_0_starting_addr strg_ub_agg_only_agg_write_addr_gen_0_starting_addr_inst0 (
    .I(config_reg_9_O),
    .O(strg_ub_agg_only_agg_write_addr_gen_0_starting_addr_inst0_O)
);
strg_ub_agg_only_agg_write_addr_gen_0_strides_0 strg_ub_agg_only_agg_write_addr_gen_0_strides_0_inst0 (
    .I(config_reg_9_O),
    .O(strg_ub_agg_only_agg_write_addr_gen_0_strides_0_inst0_O)
);
strg_ub_agg_only_agg_write_addr_gen_0_strides_1 strg_ub_agg_only_agg_write_addr_gen_0_strides_1_inst0 (
    .I(config_reg_10_O),
    .O(strg_ub_agg_only_agg_write_addr_gen_0_strides_1_inst0_O)
);
strg_ub_agg_only_agg_write_addr_gen_0_strides_2 strg_ub_agg_only_agg_write_addr_gen_0_strides_2_inst0 (
    .I(config_reg_10_O),
    .O(strg_ub_agg_only_agg_write_addr_gen_0_strides_2_inst0_O)
);
strg_ub_agg_only_agg_write_addr_gen_0_strides_3 strg_ub_agg_only_agg_write_addr_gen_0_strides_3_inst0 (
    .I(config_reg_10_O),
    .O(strg_ub_agg_only_agg_write_addr_gen_0_strides_3_inst0_O)
);
strg_ub_agg_only_agg_write_addr_gen_0_strides_4 strg_ub_agg_only_agg_write_addr_gen_0_strides_4_inst0 (
    .I(config_reg_10_O),
    .O(strg_ub_agg_only_agg_write_addr_gen_0_strides_4_inst0_O)
);
strg_ub_agg_only_agg_write_addr_gen_0_strides_5 strg_ub_agg_only_agg_write_addr_gen_0_strides_5_inst0 (
    .I(config_reg_10_O),
    .O(strg_ub_agg_only_agg_write_addr_gen_0_strides_5_inst0_O)
);
strg_ub_agg_only_agg_write_addr_gen_1_starting_addr strg_ub_agg_only_agg_write_addr_gen_1_starting_addr_inst0 (
    .I(config_reg_10_O),
    .O(strg_ub_agg_only_agg_write_addr_gen_1_starting_addr_inst0_O)
);
strg_ub_agg_only_agg_write_addr_gen_1_strides_0 strg_ub_agg_only_agg_write_addr_gen_1_strides_0_inst0 (
    .I(config_reg_10_O),
    .O(strg_ub_agg_only_agg_write_addr_gen_1_strides_0_inst0_O)
);
strg_ub_agg_only_agg_write_addr_gen_1_strides_1 strg_ub_agg_only_agg_write_addr_gen_1_strides_1_inst0 (
    .I(config_reg_10_O),
    .O(strg_ub_agg_only_agg_write_addr_gen_1_strides_1_inst0_O)
);
strg_ub_agg_only_agg_write_addr_gen_1_strides_2 strg_ub_agg_only_agg_write_addr_gen_1_strides_2_inst0 (
    .I(config_reg_11_O),
    .O(strg_ub_agg_only_agg_write_addr_gen_1_strides_2_inst0_O)
);
strg_ub_agg_only_agg_write_addr_gen_1_strides_3 strg_ub_agg_only_agg_write_addr_gen_1_strides_3_inst0 (
    .I(config_reg_11_O),
    .O(strg_ub_agg_only_agg_write_addr_gen_1_strides_3_inst0_O)
);
strg_ub_agg_only_agg_write_addr_gen_1_strides_4 strg_ub_agg_only_agg_write_addr_gen_1_strides_4_inst0 (
    .I(config_reg_11_O),
    .O(strg_ub_agg_only_agg_write_addr_gen_1_strides_4_inst0_O)
);
strg_ub_agg_only_agg_write_addr_gen_1_strides_5 strg_ub_agg_only_agg_write_addr_gen_1_strides_5_inst0 (
    .I(config_reg_11_O),
    .O(strg_ub_agg_only_agg_write_addr_gen_1_strides_5_inst0_O)
);
strg_ub_agg_only_agg_write_sched_gen_0_enable strg_ub_agg_only_agg_write_sched_gen_0_enable_inst0 (
    .I(config_reg_11_O),
    .O(strg_ub_agg_only_agg_write_sched_gen_0_enable_inst0_O)
);
strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr_inst0 (
    .I(config_reg_12_O),
    .O(strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_starting_addr_inst0_O)
);
strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0 strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0_inst0 (
    .I(config_reg_12_O),
    .O(strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_0_inst0_O)
);
strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1 strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1_inst0 (
    .I(config_reg_13_O),
    .O(strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_1_inst0_O)
);
strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2 strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2_inst0 (
    .I(config_reg_13_O),
    .O(strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_2_inst0_O)
);
strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3 strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3_inst0 (
    .I(config_reg_14_O),
    .O(strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_3_inst0_O)
);
strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4 strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4_inst0 (
    .I(config_reg_14_O),
    .O(strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_4_inst0_O)
);
strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5 strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5_inst0 (
    .I(config_reg_15_O),
    .O(strg_ub_agg_only_agg_write_sched_gen_0_sched_addr_gen_strides_5_inst0_O)
);
strg_ub_agg_only_agg_write_sched_gen_1_enable strg_ub_agg_only_agg_write_sched_gen_1_enable_inst0 (
    .I(config_reg_15_O),
    .O(strg_ub_agg_only_agg_write_sched_gen_1_enable_inst0_O)
);
strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr_inst0 (
    .I(config_reg_16_O),
    .O(strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_starting_addr_inst0_O)
);
strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0 strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0_inst0 (
    .I(config_reg_16_O),
    .O(strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_0_inst0_O)
);
strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1 strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1_inst0 (
    .I(config_reg_17_O),
    .O(strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_1_inst0_O)
);
strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2 strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2_inst0 (
    .I(config_reg_17_O),
    .O(strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_2_inst0_O)
);
strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3 strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3_inst0 (
    .I(config_reg_18_O),
    .O(strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_3_inst0_O)
);
strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4 strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4_inst0 (
    .I(config_reg_18_O),
    .O(strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_4_inst0_O)
);
strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5 strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5_inst0 (
    .I(config_reg_19_O),
    .O(strg_ub_agg_only_agg_write_sched_gen_1_sched_addr_gen_strides_5_inst0_O)
);
strg_ub_agg_only_loops_in2buf_0_dimensionality strg_ub_agg_only_loops_in2buf_0_dimensionality_inst0 (
    .I(config_reg_19_O),
    .O(strg_ub_agg_only_loops_in2buf_0_dimensionality_inst0_O)
);
strg_ub_agg_only_loops_in2buf_0_ranges_0 strg_ub_agg_only_loops_in2buf_0_ranges_0_inst0 (
    .I(config_reg_20_O),
    .O(strg_ub_agg_only_loops_in2buf_0_ranges_0_inst0_O)
);
strg_ub_agg_only_loops_in2buf_0_ranges_1 strg_ub_agg_only_loops_in2buf_0_ranges_1_inst0 (
    .I(config_reg_20_O),
    .O(strg_ub_agg_only_loops_in2buf_0_ranges_1_inst0_O)
);
strg_ub_agg_only_loops_in2buf_0_ranges_2 strg_ub_agg_only_loops_in2buf_0_ranges_2_inst0 (
    .I(config_reg_21_O),
    .O(strg_ub_agg_only_loops_in2buf_0_ranges_2_inst0_O)
);
strg_ub_agg_only_loops_in2buf_0_ranges_3 strg_ub_agg_only_loops_in2buf_0_ranges_3_inst0 (
    .I(config_reg_21_O),
    .O(strg_ub_agg_only_loops_in2buf_0_ranges_3_inst0_O)
);
strg_ub_agg_only_loops_in2buf_0_ranges_4 strg_ub_agg_only_loops_in2buf_0_ranges_4_inst0 (
    .I(config_reg_22_O),
    .O(strg_ub_agg_only_loops_in2buf_0_ranges_4_inst0_O)
);
strg_ub_agg_only_loops_in2buf_0_ranges_5 strg_ub_agg_only_loops_in2buf_0_ranges_5_inst0 (
    .I(config_reg_22_O),
    .O(strg_ub_agg_only_loops_in2buf_0_ranges_5_inst0_O)
);
strg_ub_agg_only_loops_in2buf_1_dimensionality strg_ub_agg_only_loops_in2buf_1_dimensionality_inst0 (
    .I(config_reg_23_O),
    .O(strg_ub_agg_only_loops_in2buf_1_dimensionality_inst0_O)
);
strg_ub_agg_only_loops_in2buf_1_ranges_0 strg_ub_agg_only_loops_in2buf_1_ranges_0_inst0 (
    .I(config_reg_23_O),
    .O(strg_ub_agg_only_loops_in2buf_1_ranges_0_inst0_O)
);
strg_ub_agg_only_loops_in2buf_1_ranges_1 strg_ub_agg_only_loops_in2buf_1_ranges_1_inst0 (
    .I(config_reg_24_O),
    .O(strg_ub_agg_only_loops_in2buf_1_ranges_1_inst0_O)
);
strg_ub_agg_only_loops_in2buf_1_ranges_2 strg_ub_agg_only_loops_in2buf_1_ranges_2_inst0 (
    .I(config_reg_24_O),
    .O(strg_ub_agg_only_loops_in2buf_1_ranges_2_inst0_O)
);
strg_ub_agg_only_loops_in2buf_1_ranges_3 strg_ub_agg_only_loops_in2buf_1_ranges_3_inst0 (
    .I(config_reg_25_O),
    .O(strg_ub_agg_only_loops_in2buf_1_ranges_3_inst0_O)
);
strg_ub_agg_only_loops_in2buf_1_ranges_4 strg_ub_agg_only_loops_in2buf_1_ranges_4_inst0 (
    .I(config_reg_25_O),
    .O(strg_ub_agg_only_loops_in2buf_1_ranges_4_inst0_O)
);
strg_ub_agg_only_loops_in2buf_1_ranges_5 strg_ub_agg_only_loops_in2buf_1_ranges_5_inst0 (
    .I(config_reg_26_O),
    .O(strg_ub_agg_only_loops_in2buf_1_ranges_5_inst0_O)
);
strg_ub_agg_sram_shared_agg_read_sched_gen_0_enable strg_ub_agg_sram_shared_agg_read_sched_gen_0_enable_inst0 (
    .I(config_reg_26_O),
    .O(strg_ub_agg_sram_shared_agg_read_sched_gen_0_enable_inst0_O)
);
strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr_inst0 (
    .I(config_reg_27_O),
    .O(strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_starting_addr_inst0_O)
);
strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0 strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0_inst0 (
    .I(config_reg_27_O),
    .O(strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_0_inst0_O)
);
strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1 strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1_inst0 (
    .I(config_reg_28_O),
    .O(strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_1_inst0_O)
);
strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2 strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2_inst0 (
    .I(config_reg_28_O),
    .O(strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_2_inst0_O)
);
strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3 strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3_inst0 (
    .I(config_reg_29_O),
    .O(strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_3_inst0_O)
);
strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4 strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4_inst0 (
    .I(config_reg_29_O),
    .O(strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_4_inst0_O)
);
strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5 strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5_inst0 (
    .I(config_reg_30_O),
    .O(strg_ub_agg_sram_shared_agg_read_sched_gen_0_sched_addr_gen_strides_5_inst0_O)
);
strg_ub_agg_sram_shared_agg_read_sched_gen_1_enable strg_ub_agg_sram_shared_agg_read_sched_gen_1_enable_inst0 (
    .I(config_reg_30_O),
    .O(strg_ub_agg_sram_shared_agg_read_sched_gen_1_enable_inst0_O)
);
strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr_inst0 (
    .I(config_reg_31_O),
    .O(strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_starting_addr_inst0_O)
);
strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0 strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0_inst0 (
    .I(config_reg_31_O),
    .O(strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_0_inst0_O)
);
strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1 strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1_inst0 (
    .I(config_reg_32_O),
    .O(strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_1_inst0_O)
);
strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2 strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2_inst0 (
    .I(config_reg_32_O),
    .O(strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_2_inst0_O)
);
strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3 strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3_inst0 (
    .I(config_reg_33_O),
    .O(strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_3_inst0_O)
);
strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4 strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4_inst0 (
    .I(config_reg_33_O),
    .O(strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_4_inst0_O)
);
strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5 strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5_inst0 (
    .I(config_reg_34_O),
    .O(strg_ub_agg_sram_shared_agg_read_sched_gen_1_sched_addr_gen_strides_5_inst0_O)
);
strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality_inst0 (
    .I(config_reg_34_O),
    .O(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_dimensionality_inst0_O)
);
strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0 strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0_inst0 (
    .I(config_reg_35_O),
    .O(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_0_inst0_O)
);
strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1 strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1_inst0 (
    .I(config_reg_35_O),
    .O(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_1_inst0_O)
);
strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2 strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2_inst0 (
    .I(config_reg_36_O),
    .O(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_2_inst0_O)
);
strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3 strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3_inst0 (
    .I(config_reg_36_O),
    .O(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_3_inst0_O)
);
strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4 strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4_inst0 (
    .I(config_reg_37_O),
    .O(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_4_inst0_O)
);
strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5 strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5_inst0 (
    .I(config_reg_37_O),
    .O(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_0_ranges_5_inst0_O)
);
strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality_inst0 (
    .I(config_reg_38_O),
    .O(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_dimensionality_inst0_O)
);
strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0 strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0_inst0 (
    .I(config_reg_38_O),
    .O(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_0_inst0_O)
);
strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1 strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1_inst0 (
    .I(config_reg_39_O),
    .O(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_1_inst0_O)
);
strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2 strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2_inst0 (
    .I(config_reg_39_O),
    .O(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_2_inst0_O)
);
strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3 strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3_inst0 (
    .I(config_reg_40_O),
    .O(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_3_inst0_O)
);
strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4 strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4_inst0 (
    .I(config_reg_40_O),
    .O(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_4_inst0_O)
);
strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5 strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5_inst0 (
    .I(config_reg_41_O),
    .O(strg_ub_agg_sram_shared_loops_in2buf_autovec_write_1_ranges_5_inst0_O)
);
strg_ub_sram_only_input_addr_gen_0_starting_addr strg_ub_sram_only_input_addr_gen_0_starting_addr_inst0 (
    .I(config_reg_41_O),
    .O(strg_ub_sram_only_input_addr_gen_0_starting_addr_inst0_O)
);
strg_ub_sram_only_input_addr_gen_0_strides_0 strg_ub_sram_only_input_addr_gen_0_strides_0_inst0 (
    .I(config_reg_42_O),
    .O(strg_ub_sram_only_input_addr_gen_0_strides_0_inst0_O)
);
strg_ub_sram_only_input_addr_gen_0_strides_1 strg_ub_sram_only_input_addr_gen_0_strides_1_inst0 (
    .I(config_reg_42_O),
    .O(strg_ub_sram_only_input_addr_gen_0_strides_1_inst0_O)
);
strg_ub_sram_only_input_addr_gen_0_strides_2 strg_ub_sram_only_input_addr_gen_0_strides_2_inst0 (
    .I(config_reg_42_O),
    .O(strg_ub_sram_only_input_addr_gen_0_strides_2_inst0_O)
);
strg_ub_sram_only_input_addr_gen_0_strides_3 strg_ub_sram_only_input_addr_gen_0_strides_3_inst0 (
    .I(config_reg_43_O),
    .O(strg_ub_sram_only_input_addr_gen_0_strides_3_inst0_O)
);
strg_ub_sram_only_input_addr_gen_0_strides_4 strg_ub_sram_only_input_addr_gen_0_strides_4_inst0 (
    .I(config_reg_43_O),
    .O(strg_ub_sram_only_input_addr_gen_0_strides_4_inst0_O)
);
strg_ub_sram_only_input_addr_gen_0_strides_5 strg_ub_sram_only_input_addr_gen_0_strides_5_inst0 (
    .I(config_reg_43_O),
    .O(strg_ub_sram_only_input_addr_gen_0_strides_5_inst0_O)
);
strg_ub_sram_only_input_addr_gen_1_starting_addr strg_ub_sram_only_input_addr_gen_1_starting_addr_inst0 (
    .I(config_reg_44_O),
    .O(strg_ub_sram_only_input_addr_gen_1_starting_addr_inst0_O)
);
strg_ub_sram_only_input_addr_gen_1_strides_0 strg_ub_sram_only_input_addr_gen_1_strides_0_inst0 (
    .I(config_reg_44_O),
    .O(strg_ub_sram_only_input_addr_gen_1_strides_0_inst0_O)
);
strg_ub_sram_only_input_addr_gen_1_strides_1 strg_ub_sram_only_input_addr_gen_1_strides_1_inst0 (
    .I(config_reg_44_O),
    .O(strg_ub_sram_only_input_addr_gen_1_strides_1_inst0_O)
);
strg_ub_sram_only_input_addr_gen_1_strides_2 strg_ub_sram_only_input_addr_gen_1_strides_2_inst0 (
    .I(config_reg_45_O),
    .O(strg_ub_sram_only_input_addr_gen_1_strides_2_inst0_O)
);
strg_ub_sram_only_input_addr_gen_1_strides_3 strg_ub_sram_only_input_addr_gen_1_strides_3_inst0 (
    .I(config_reg_45_O),
    .O(strg_ub_sram_only_input_addr_gen_1_strides_3_inst0_O)
);
strg_ub_sram_only_input_addr_gen_1_strides_4 strg_ub_sram_only_input_addr_gen_1_strides_4_inst0 (
    .I(config_reg_45_O),
    .O(strg_ub_sram_only_input_addr_gen_1_strides_4_inst0_O)
);
strg_ub_sram_only_input_addr_gen_1_strides_5 strg_ub_sram_only_input_addr_gen_1_strides_5_inst0 (
    .I(config_reg_46_O),
    .O(strg_ub_sram_only_input_addr_gen_1_strides_5_inst0_O)
);
strg_ub_sram_only_output_addr_gen_0_starting_addr strg_ub_sram_only_output_addr_gen_0_starting_addr_inst0 (
    .I(config_reg_46_O),
    .O(strg_ub_sram_only_output_addr_gen_0_starting_addr_inst0_O)
);
strg_ub_sram_only_output_addr_gen_0_strides_0 strg_ub_sram_only_output_addr_gen_0_strides_0_inst0 (
    .I(config_reg_46_O),
    .O(strg_ub_sram_only_output_addr_gen_0_strides_0_inst0_O)
);
strg_ub_sram_only_output_addr_gen_0_strides_1 strg_ub_sram_only_output_addr_gen_0_strides_1_inst0 (
    .I(config_reg_47_O),
    .O(strg_ub_sram_only_output_addr_gen_0_strides_1_inst0_O)
);
strg_ub_sram_only_output_addr_gen_0_strides_2 strg_ub_sram_only_output_addr_gen_0_strides_2_inst0 (
    .I(config_reg_47_O),
    .O(strg_ub_sram_only_output_addr_gen_0_strides_2_inst0_O)
);
strg_ub_sram_only_output_addr_gen_0_strides_3 strg_ub_sram_only_output_addr_gen_0_strides_3_inst0 (
    .I(config_reg_47_O),
    .O(strg_ub_sram_only_output_addr_gen_0_strides_3_inst0_O)
);
strg_ub_sram_only_output_addr_gen_0_strides_4 strg_ub_sram_only_output_addr_gen_0_strides_4_inst0 (
    .I(config_reg_48_O),
    .O(strg_ub_sram_only_output_addr_gen_0_strides_4_inst0_O)
);
strg_ub_sram_only_output_addr_gen_0_strides_5 strg_ub_sram_only_output_addr_gen_0_strides_5_inst0 (
    .I(config_reg_48_O),
    .O(strg_ub_sram_only_output_addr_gen_0_strides_5_inst0_O)
);
strg_ub_sram_only_output_addr_gen_1_starting_addr strg_ub_sram_only_output_addr_gen_1_starting_addr_inst0 (
    .I(config_reg_48_O),
    .O(strg_ub_sram_only_output_addr_gen_1_starting_addr_inst0_O)
);
strg_ub_sram_only_output_addr_gen_1_strides_0 strg_ub_sram_only_output_addr_gen_1_strides_0_inst0 (
    .I(config_reg_49_O),
    .O(strg_ub_sram_only_output_addr_gen_1_strides_0_inst0_O)
);
strg_ub_sram_only_output_addr_gen_1_strides_1 strg_ub_sram_only_output_addr_gen_1_strides_1_inst0 (
    .I(config_reg_49_O),
    .O(strg_ub_sram_only_output_addr_gen_1_strides_1_inst0_O)
);
strg_ub_sram_only_output_addr_gen_1_strides_2 strg_ub_sram_only_output_addr_gen_1_strides_2_inst0 (
    .I(config_reg_49_O),
    .O(strg_ub_sram_only_output_addr_gen_1_strides_2_inst0_O)
);
strg_ub_sram_only_output_addr_gen_1_strides_3 strg_ub_sram_only_output_addr_gen_1_strides_3_inst0 (
    .I(config_reg_50_O),
    .O(strg_ub_sram_only_output_addr_gen_1_strides_3_inst0_O)
);
strg_ub_sram_only_output_addr_gen_1_strides_4 strg_ub_sram_only_output_addr_gen_1_strides_4_inst0 (
    .I(config_reg_50_O),
    .O(strg_ub_sram_only_output_addr_gen_1_strides_4_inst0_O)
);
strg_ub_sram_only_output_addr_gen_1_strides_5 strg_ub_sram_only_output_addr_gen_1_strides_5_inst0 (
    .I(config_reg_50_O),
    .O(strg_ub_sram_only_output_addr_gen_1_strides_5_inst0_O)
);
strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality_inst0 (
    .I(config_reg_50_O),
    .O(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_dimensionality_inst0_O)
);
strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0 strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0_inst0 (
    .I(config_reg_51_O),
    .O(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_0_inst0_O)
);
strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1 strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1_inst0 (
    .I(config_reg_51_O),
    .O(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_1_inst0_O)
);
strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2 strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2_inst0 (
    .I(config_reg_52_O),
    .O(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_2_inst0_O)
);
strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3 strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3_inst0 (
    .I(config_reg_52_O),
    .O(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_3_inst0_O)
);
strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4 strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4_inst0 (
    .I(config_reg_53_O),
    .O(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_4_inst0_O)
);
strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5 strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5_inst0 (
    .I(config_reg_53_O),
    .O(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_0_ranges_5_inst0_O)
);
strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality_inst0 (
    .I(config_reg_54_O),
    .O(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_dimensionality_inst0_O)
);
strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0 strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0_inst0 (
    .I(config_reg_54_O),
    .O(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_0_inst0_O)
);
strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1 strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1_inst0 (
    .I(config_reg_55_O),
    .O(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_1_inst0_O)
);
strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2 strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2_inst0 (
    .I(config_reg_55_O),
    .O(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_2_inst0_O)
);
strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3 strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3_inst0 (
    .I(config_reg_56_O),
    .O(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_3_inst0_O)
);
strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4 strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4_inst0 (
    .I(config_reg_56_O),
    .O(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_4_inst0_O)
);
strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5 strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5_inst0 (
    .I(config_reg_57_O),
    .O(strg_ub_sram_tb_shared_loops_buf2out_autovec_read_1_ranges_5_inst0_O)
);
strg_ub_sram_tb_shared_output_sched_gen_0_enable strg_ub_sram_tb_shared_output_sched_gen_0_enable_inst0 (
    .I(config_reg_57_O),
    .O(strg_ub_sram_tb_shared_output_sched_gen_0_enable_inst0_O)
);
strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr_inst0 (
    .I(config_reg_58_O),
    .O(strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_starting_addr_inst0_O)
);
strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0 strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0_inst0 (
    .I(config_reg_58_O),
    .O(strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_0_inst0_O)
);
strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1 strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1_inst0 (
    .I(config_reg_59_O),
    .O(strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_1_inst0_O)
);
strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2 strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2_inst0 (
    .I(config_reg_59_O),
    .O(strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_2_inst0_O)
);
strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3 strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3_inst0 (
    .I(config_reg_60_O),
    .O(strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_3_inst0_O)
);
strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4 strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4_inst0 (
    .I(config_reg_60_O),
    .O(strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_4_inst0_O)
);
strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5 strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5_inst0 (
    .I(config_reg_61_O),
    .O(strg_ub_sram_tb_shared_output_sched_gen_0_sched_addr_gen_strides_5_inst0_O)
);
strg_ub_sram_tb_shared_output_sched_gen_1_enable strg_ub_sram_tb_shared_output_sched_gen_1_enable_inst0 (
    .I(config_reg_61_O),
    .O(strg_ub_sram_tb_shared_output_sched_gen_1_enable_inst0_O)
);
strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr_inst0 (
    .I(config_reg_62_O),
    .O(strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_starting_addr_inst0_O)
);
strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0 strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0_inst0 (
    .I(config_reg_62_O),
    .O(strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_0_inst0_O)
);
strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1 strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1_inst0 (
    .I(config_reg_63_O),
    .O(strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_1_inst0_O)
);
strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2 strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2_inst0 (
    .I(config_reg_63_O),
    .O(strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_2_inst0_O)
);
strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3 strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3_inst0 (
    .I(config_reg_64_O),
    .O(strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_3_inst0_O)
);
strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4 strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4_inst0 (
    .I(config_reg_64_O),
    .O(strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_4_inst0_O)
);
strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5 strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5_inst0 (
    .I(config_reg_65_O),
    .O(strg_ub_sram_tb_shared_output_sched_gen_1_sched_addr_gen_strides_5_inst0_O)
);
strg_ub_tb_only_loops_buf2out_read_0_dimensionality strg_ub_tb_only_loops_buf2out_read_0_dimensionality_inst0 (
    .I(config_reg_65_O),
    .O(strg_ub_tb_only_loops_buf2out_read_0_dimensionality_inst0_O)
);
strg_ub_tb_only_loops_buf2out_read_0_ranges_0 strg_ub_tb_only_loops_buf2out_read_0_ranges_0_inst0 (
    .I(config_reg_66_O),
    .O(strg_ub_tb_only_loops_buf2out_read_0_ranges_0_inst0_O)
);
strg_ub_tb_only_loops_buf2out_read_0_ranges_1 strg_ub_tb_only_loops_buf2out_read_0_ranges_1_inst0 (
    .I(config_reg_66_O),
    .O(strg_ub_tb_only_loops_buf2out_read_0_ranges_1_inst0_O)
);
strg_ub_tb_only_loops_buf2out_read_0_ranges_2 strg_ub_tb_only_loops_buf2out_read_0_ranges_2_inst0 (
    .I(config_reg_67_O),
    .O(strg_ub_tb_only_loops_buf2out_read_0_ranges_2_inst0_O)
);
strg_ub_tb_only_loops_buf2out_read_0_ranges_3 strg_ub_tb_only_loops_buf2out_read_0_ranges_3_inst0 (
    .I(config_reg_67_O),
    .O(strg_ub_tb_only_loops_buf2out_read_0_ranges_3_inst0_O)
);
strg_ub_tb_only_loops_buf2out_read_0_ranges_4 strg_ub_tb_only_loops_buf2out_read_0_ranges_4_inst0 (
    .I(config_reg_68_O),
    .O(strg_ub_tb_only_loops_buf2out_read_0_ranges_4_inst0_O)
);
strg_ub_tb_only_loops_buf2out_read_0_ranges_5 strg_ub_tb_only_loops_buf2out_read_0_ranges_5_inst0 (
    .I(config_reg_68_O),
    .O(strg_ub_tb_only_loops_buf2out_read_0_ranges_5_inst0_O)
);
strg_ub_tb_only_loops_buf2out_read_1_dimensionality strg_ub_tb_only_loops_buf2out_read_1_dimensionality_inst0 (
    .I(config_reg_69_O),
    .O(strg_ub_tb_only_loops_buf2out_read_1_dimensionality_inst0_O)
);
strg_ub_tb_only_loops_buf2out_read_1_ranges_0 strg_ub_tb_only_loops_buf2out_read_1_ranges_0_inst0 (
    .I(config_reg_69_O),
    .O(strg_ub_tb_only_loops_buf2out_read_1_ranges_0_inst0_O)
);
strg_ub_tb_only_loops_buf2out_read_1_ranges_1 strg_ub_tb_only_loops_buf2out_read_1_ranges_1_inst0 (
    .I(config_reg_70_O),
    .O(strg_ub_tb_only_loops_buf2out_read_1_ranges_1_inst0_O)
);
strg_ub_tb_only_loops_buf2out_read_1_ranges_2 strg_ub_tb_only_loops_buf2out_read_1_ranges_2_inst0 (
    .I(config_reg_70_O),
    .O(strg_ub_tb_only_loops_buf2out_read_1_ranges_2_inst0_O)
);
strg_ub_tb_only_loops_buf2out_read_1_ranges_3 strg_ub_tb_only_loops_buf2out_read_1_ranges_3_inst0 (
    .I(config_reg_71_O),
    .O(strg_ub_tb_only_loops_buf2out_read_1_ranges_3_inst0_O)
);
strg_ub_tb_only_loops_buf2out_read_1_ranges_4 strg_ub_tb_only_loops_buf2out_read_1_ranges_4_inst0 (
    .I(config_reg_71_O),
    .O(strg_ub_tb_only_loops_buf2out_read_1_ranges_4_inst0_O)
);
strg_ub_tb_only_loops_buf2out_read_1_ranges_5 strg_ub_tb_only_loops_buf2out_read_1_ranges_5_inst0 (
    .I(config_reg_72_O),
    .O(strg_ub_tb_only_loops_buf2out_read_1_ranges_5_inst0_O)
);
strg_ub_tb_only_tb_read_addr_gen_0_starting_addr strg_ub_tb_only_tb_read_addr_gen_0_starting_addr_inst0 (
    .I(config_reg_72_O),
    .O(strg_ub_tb_only_tb_read_addr_gen_0_starting_addr_inst0_O)
);
strg_ub_tb_only_tb_read_addr_gen_0_strides_0 strg_ub_tb_only_tb_read_addr_gen_0_strides_0_inst0 (
    .I(config_reg_72_O),
    .O(strg_ub_tb_only_tb_read_addr_gen_0_strides_0_inst0_O)
);
strg_ub_tb_only_tb_read_addr_gen_0_strides_1 strg_ub_tb_only_tb_read_addr_gen_0_strides_1_inst0 (
    .I(config_reg_72_O),
    .O(strg_ub_tb_only_tb_read_addr_gen_0_strides_1_inst0_O)
);
strg_ub_tb_only_tb_read_addr_gen_0_strides_2 strg_ub_tb_only_tb_read_addr_gen_0_strides_2_inst0 (
    .I(config_reg_72_O),
    .O(strg_ub_tb_only_tb_read_addr_gen_0_strides_2_inst0_O)
);
strg_ub_tb_only_tb_read_addr_gen_0_strides_3 strg_ub_tb_only_tb_read_addr_gen_0_strides_3_inst0 (
    .I(config_reg_73_O),
    .O(strg_ub_tb_only_tb_read_addr_gen_0_strides_3_inst0_O)
);
strg_ub_tb_only_tb_read_addr_gen_0_strides_4 strg_ub_tb_only_tb_read_addr_gen_0_strides_4_inst0 (
    .I(config_reg_73_O),
    .O(strg_ub_tb_only_tb_read_addr_gen_0_strides_4_inst0_O)
);
strg_ub_tb_only_tb_read_addr_gen_0_strides_5 strg_ub_tb_only_tb_read_addr_gen_0_strides_5_inst0 (
    .I(config_reg_73_O),
    .O(strg_ub_tb_only_tb_read_addr_gen_0_strides_5_inst0_O)
);
strg_ub_tb_only_tb_read_addr_gen_1_starting_addr strg_ub_tb_only_tb_read_addr_gen_1_starting_addr_inst0 (
    .I(config_reg_73_O),
    .O(strg_ub_tb_only_tb_read_addr_gen_1_starting_addr_inst0_O)
);
strg_ub_tb_only_tb_read_addr_gen_1_strides_0 strg_ub_tb_only_tb_read_addr_gen_1_strides_0_inst0 (
    .I(config_reg_73_O),
    .O(strg_ub_tb_only_tb_read_addr_gen_1_strides_0_inst0_O)
);
strg_ub_tb_only_tb_read_addr_gen_1_strides_1 strg_ub_tb_only_tb_read_addr_gen_1_strides_1_inst0 (
    .I(config_reg_73_O),
    .O(strg_ub_tb_only_tb_read_addr_gen_1_strides_1_inst0_O)
);
strg_ub_tb_only_tb_read_addr_gen_1_strides_2 strg_ub_tb_only_tb_read_addr_gen_1_strides_2_inst0 (
    .I(config_reg_73_O),
    .O(strg_ub_tb_only_tb_read_addr_gen_1_strides_2_inst0_O)
);
strg_ub_tb_only_tb_read_addr_gen_1_strides_3 strg_ub_tb_only_tb_read_addr_gen_1_strides_3_inst0 (
    .I(config_reg_73_O),
    .O(strg_ub_tb_only_tb_read_addr_gen_1_strides_3_inst0_O)
);
strg_ub_tb_only_tb_read_addr_gen_1_strides_4 strg_ub_tb_only_tb_read_addr_gen_1_strides_4_inst0 (
    .I(config_reg_74_O),
    .O(strg_ub_tb_only_tb_read_addr_gen_1_strides_4_inst0_O)
);
strg_ub_tb_only_tb_read_addr_gen_1_strides_5 strg_ub_tb_only_tb_read_addr_gen_1_strides_5_inst0 (
    .I(config_reg_74_O),
    .O(strg_ub_tb_only_tb_read_addr_gen_1_strides_5_inst0_O)
);
strg_ub_tb_only_tb_read_sched_gen_0_enable strg_ub_tb_only_tb_read_sched_gen_0_enable_inst0 (
    .I(config_reg_74_O),
    .O(strg_ub_tb_only_tb_read_sched_gen_0_enable_inst0_O)
);
strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr_inst0 (
    .I(config_reg_74_O),
    .O(strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_starting_addr_inst0_O)
);
strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0 strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0_inst0 (
    .I(config_reg_75_O),
    .O(strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_0_inst0_O)
);
strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1 strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1_inst0 (
    .I(config_reg_75_O),
    .O(strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_1_inst0_O)
);
strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2 strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2_inst0 (
    .I(config_reg_76_O),
    .O(strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_2_inst0_O)
);
strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3 strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3_inst0 (
    .I(config_reg_76_O),
    .O(strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_3_inst0_O)
);
strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4 strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4_inst0 (
    .I(config_reg_77_O),
    .O(strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_4_inst0_O)
);
strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5 strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5_inst0 (
    .I(config_reg_77_O),
    .O(strg_ub_tb_only_tb_read_sched_gen_0_sched_addr_gen_strides_5_inst0_O)
);
strg_ub_tb_only_tb_read_sched_gen_1_enable strg_ub_tb_only_tb_read_sched_gen_1_enable_inst0 (
    .I(config_reg_78_O),
    .O(strg_ub_tb_only_tb_read_sched_gen_1_enable_inst0_O)
);
strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr_inst0 (
    .I(config_reg_78_O),
    .O(strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_starting_addr_inst0_O)
);
strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0 strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0_inst0 (
    .I(config_reg_79_O),
    .O(strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_0_inst0_O)
);
strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1 strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1_inst0 (
    .I(config_reg_79_O),
    .O(strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_1_inst0_O)
);
strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2 strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2_inst0 (
    .I(config_reg_80_O),
    .O(strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_2_inst0_O)
);
strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3 strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3_inst0 (
    .I(config_reg_80_O),
    .O(strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_3_inst0_O)
);
strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4 strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4_inst0 (
    .I(config_reg_81_O),
    .O(strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_4_inst0_O)
);
strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5 strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5_inst0 (
    .I(config_reg_81_O),
    .O(strg_ub_tb_only_tb_read_sched_gen_1_sched_addr_gen_strides_5_inst0_O)
);
strg_ub_tb_only_tb_write_addr_gen_0_starting_addr strg_ub_tb_only_tb_write_addr_gen_0_starting_addr_inst0 (
    .I(config_reg_82_O),
    .O(strg_ub_tb_only_tb_write_addr_gen_0_starting_addr_inst0_O)
);
strg_ub_tb_only_tb_write_addr_gen_0_strides_0 strg_ub_tb_only_tb_write_addr_gen_0_strides_0_inst0 (
    .I(config_reg_82_O),
    .O(strg_ub_tb_only_tb_write_addr_gen_0_strides_0_inst0_O)
);
strg_ub_tb_only_tb_write_addr_gen_0_strides_1 strg_ub_tb_only_tb_write_addr_gen_0_strides_1_inst0 (
    .I(config_reg_82_O),
    .O(strg_ub_tb_only_tb_write_addr_gen_0_strides_1_inst0_O)
);
strg_ub_tb_only_tb_write_addr_gen_0_strides_2 strg_ub_tb_only_tb_write_addr_gen_0_strides_2_inst0 (
    .I(config_reg_82_O),
    .O(strg_ub_tb_only_tb_write_addr_gen_0_strides_2_inst0_O)
);
strg_ub_tb_only_tb_write_addr_gen_0_strides_3 strg_ub_tb_only_tb_write_addr_gen_0_strides_3_inst0 (
    .I(config_reg_82_O),
    .O(strg_ub_tb_only_tb_write_addr_gen_0_strides_3_inst0_O)
);
strg_ub_tb_only_tb_write_addr_gen_0_strides_4 strg_ub_tb_only_tb_write_addr_gen_0_strides_4_inst0 (
    .I(config_reg_82_O),
    .O(strg_ub_tb_only_tb_write_addr_gen_0_strides_4_inst0_O)
);
strg_ub_tb_only_tb_write_addr_gen_0_strides_5 strg_ub_tb_only_tb_write_addr_gen_0_strides_5_inst0 (
    .I(config_reg_82_O),
    .O(strg_ub_tb_only_tb_write_addr_gen_0_strides_5_inst0_O)
);
strg_ub_tb_only_tb_write_addr_gen_1_starting_addr strg_ub_tb_only_tb_write_addr_gen_1_starting_addr_inst0 (
    .I(config_reg_82_O),
    .O(strg_ub_tb_only_tb_write_addr_gen_1_starting_addr_inst0_O)
);
strg_ub_tb_only_tb_write_addr_gen_1_strides_0 strg_ub_tb_only_tb_write_addr_gen_1_strides_0_inst0 (
    .I(config_reg_83_O),
    .O(strg_ub_tb_only_tb_write_addr_gen_1_strides_0_inst0_O)
);
strg_ub_tb_only_tb_write_addr_gen_1_strides_1 strg_ub_tb_only_tb_write_addr_gen_1_strides_1_inst0 (
    .I(config_reg_83_O),
    .O(strg_ub_tb_only_tb_write_addr_gen_1_strides_1_inst0_O)
);
strg_ub_tb_only_tb_write_addr_gen_1_strides_2 strg_ub_tb_only_tb_write_addr_gen_1_strides_2_inst0 (
    .I(config_reg_83_O),
    .O(strg_ub_tb_only_tb_write_addr_gen_1_strides_2_inst0_O)
);
strg_ub_tb_only_tb_write_addr_gen_1_strides_3 strg_ub_tb_only_tb_write_addr_gen_1_strides_3_inst0 (
    .I(config_reg_83_O),
    .O(strg_ub_tb_only_tb_write_addr_gen_1_strides_3_inst0_O)
);
strg_ub_tb_only_tb_write_addr_gen_1_strides_4 strg_ub_tb_only_tb_write_addr_gen_1_strides_4_inst0 (
    .I(config_reg_83_O),
    .O(strg_ub_tb_only_tb_write_addr_gen_1_strides_4_inst0_O)
);
strg_ub_tb_only_tb_write_addr_gen_1_strides_5 strg_ub_tb_only_tb_write_addr_gen_1_strides_5_inst0 (
    .I(config_reg_83_O),
    .O(strg_ub_tb_only_tb_write_addr_gen_1_strides_5_inst0_O)
);
tile_en tile_en_inst0 (
    .I(config_reg_83_O),
    .O(tile_en_inst0_O)
);
wen_in_0_reg_sel wen_in_0_reg_sel_inst0 (
    .I(config_reg_83_O),
    .O(wen_in_0_reg_sel_inst0_O)
);
wen_in_0_reg_value wen_in_0_reg_value_inst0 (
    .I(config_reg_83_O),
    .O(wen_in_0_reg_value_inst0_O)
);
coreir_mux #(
    .width(1)
) wen_in_0_sel$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(wen_in_0),
    .in1(wen_in_0_reg_value_inst0_O),
    .sel(wen_in_0_reg_sel_inst0_O[0]),
    .out(wen_in_0_sel$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
wen_in_1_reg_sel wen_in_1_reg_sel_inst0 (
    .I(config_reg_83_O),
    .O(wen_in_1_reg_sel_inst0_O)
);
wen_in_1_reg_value wen_in_1_reg_value_inst0 (
    .I(config_reg_83_O),
    .O(wen_in_1_reg_value_inst0_O)
);
coreir_mux #(
    .width(1)
) wen_in_1_sel$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(wen_in_1),
    .in1(wen_in_1_reg_value_inst0_O),
    .sel(wen_in_1_reg_sel_inst0_O[0]),
    .out(wen_in_1_sel$Mux2x1_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
assign data_out_0 = LakeTop_W_inst0_data_out_0;
assign data_out_1 = LakeTop_W_inst0_data_out_1;
assign empty = LakeTop_W_inst0_empty;
assign full = LakeTop_W_inst0_full;
assign read_config_data = MuxWrapper_84_32_inst0$Mux84x32_inst0$coreir_commonlib_mux84x32_inst0_out;
assign read_config_data_1 = LakeTop_W_inst0_config_data_out_0;
assign read_config_data_2 = LakeTop_W_inst0_config_data_out_1;
assign sram_ready_out = LakeTop_W_inst0_sram_ready_out;
assign stencil_valid = LakeTop_W_inst0_stencil_valid;
assign valid_out_0 = LakeTop_W_inst0_valid_out[0];
assign valid_out_1 = LakeTop_W_inst0_valid_out[1];
endmodule

module ConfigPipeStage (
    input clk,
    input [31:0] config_config_addr,
    input [31:0] config_config_data,
    output [31:0] config_out_config_addr,
    output [31:0] config_out_config_data,
    output [0:0] config_out_read,
    output [0:0] config_out_write,
    input [0:0] config_read,
    input [0:0] config_write
);
wire [31:0] reg_P_inst0_out;
wire [31:0] reg_P_inst1_out;
wire [0:0] reg_P_inst2_out;
wire [0:0] reg_P_inst3_out;
coreir_reg #(
    .clk_posedge(1'b1),
    .init(32'h00000000),
    .width(32)
) reg_P_inst0 (
    .clk(clk),
    .in(config_config_addr),
    .out(reg_P_inst0_out)
);
coreir_reg #(
    .clk_posedge(1'b1),
    .init(32'h00000000),
    .width(32)
) reg_P_inst1 (
    .clk(clk),
    .in(config_config_data),
    .out(reg_P_inst1_out)
);
coreir_reg #(
    .clk_posedge(1'b1),
    .init(1'h0),
    .width(1)
) reg_P_inst2 (
    .clk(clk),
    .in(config_read),
    .out(reg_P_inst2_out)
);
coreir_reg #(
    .clk_posedge(1'b1),
    .init(1'h0),
    .width(1)
) reg_P_inst3 (
    .clk(clk),
    .in(config_write),
    .out(reg_P_inst3_out)
);
assign config_out_config_addr = reg_P_inst0_out;
assign config_out_config_data = reg_P_inst1_out;
assign config_out_read = reg_P_inst2_out;
assign config_out_write = reg_P_inst3_out;
endmodule

module Cond (
    input [4:0] code,
    input alu,
    input Z,
    input N,
    input C,
    input V,
    output O,
    input CLK,
    input ASYNCRESET
);
wire [0:0] Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst13$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst14$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst15$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst16$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst17$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst9$coreir_commonlib_mux2x1_inst0$_join_out;
wire [4:0] const_0_5_out;
wire [4:0] const_10_5_out;
wire [4:0] const_11_5_out;
wire [4:0] const_12_5_out;
wire [4:0] const_13_5_out;
wire [4:0] const_14_5_out;
wire [4:0] const_15_5_out;
wire [4:0] const_16_5_out;
wire [4:0] const_17_5_out;
wire [4:0] const_1_5_out;
wire [4:0] const_2_5_out;
wire [4:0] const_3_5_out;
wire [4:0] const_4_5_out;
wire [4:0] const_5_5_out;
wire [4:0] const_6_5_out;
wire [4:0] const_7_5_out;
wire [4:0] const_8_5_out;
wire [4:0] const_9_5_out;
wire magma_Bit_and_inst0_out;
wire magma_Bit_and_inst1_out;
wire magma_Bit_and_inst2_out;
wire magma_Bit_and_inst3_out;
wire magma_Bit_not_inst0_out;
wire magma_Bit_not_inst1_out;
wire magma_Bit_not_inst10_out;
wire magma_Bit_not_inst11_out;
wire magma_Bit_not_inst12_out;
wire magma_Bit_not_inst2_out;
wire magma_Bit_not_inst3_out;
wire magma_Bit_not_inst4_out;
wire magma_Bit_not_inst5_out;
wire magma_Bit_not_inst6_out;
wire magma_Bit_not_inst7_out;
wire magma_Bit_not_inst8_out;
wire magma_Bit_not_inst9_out;
wire magma_Bit_or_inst0_out;
wire magma_Bit_or_inst1_out;
wire magma_Bit_or_inst2_out;
wire magma_Bit_or_inst3_out;
wire magma_Bit_or_inst4_out;
wire magma_Bit_or_inst5_out;
wire magma_Bit_xor_inst0_out;
wire magma_Bit_xor_inst1_out;
wire magma_Bit_xor_inst2_out;
wire magma_Bit_xor_inst3_out;
wire magma_Bits_5_eq_inst0_out;
wire magma_Bits_5_eq_inst1_out;
wire magma_Bits_5_eq_inst10_out;
wire magma_Bits_5_eq_inst11_out;
wire magma_Bits_5_eq_inst12_out;
wire magma_Bits_5_eq_inst13_out;
wire magma_Bits_5_eq_inst14_out;
wire magma_Bits_5_eq_inst15_out;
wire magma_Bits_5_eq_inst16_out;
wire magma_Bits_5_eq_inst17_out;
wire magma_Bits_5_eq_inst18_out;
wire magma_Bits_5_eq_inst19_out;
wire magma_Bits_5_eq_inst2_out;
wire magma_Bits_5_eq_inst3_out;
wire magma_Bits_5_eq_inst4_out;
wire magma_Bits_5_eq_inst5_out;
wire magma_Bits_5_eq_inst6_out;
wire magma_Bits_5_eq_inst7_out;
wire magma_Bits_5_eq_inst8_out;
wire magma_Bits_5_eq_inst9_out;
coreir_mux #(
    .width(1)
) Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(magma_Bit_and_inst3_out),
    .in1(magma_Bit_or_inst5_out),
    .sel(magma_Bits_5_eq_inst0_out),
    .out(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(magma_Bit_and_inst2_out),
    .sel(magma_Bits_5_eq_inst1_out),
    .out(Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst10$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst9$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(magma_Bit_not_inst3_out),
    .sel(magma_Bits_5_eq_inst10_out),
    .out(Mux2xBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst11$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst10$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(V),
    .sel(magma_Bits_5_eq_inst11_out),
    .out(Mux2xBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst12$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst11$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(magma_Bit_not_inst2_out),
    .sel(magma_Bits_5_eq_inst12_out),
    .out(Mux2xBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst13$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst12$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(N),
    .sel(magma_Bits_5_eq_inst13_out),
    .out(Mux2xBit_inst13$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst14$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst13$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(magma_Bit_not_inst1_out),
    .sel(magma_Bit_or_inst0_out),
    .out(Mux2xBit_inst14$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst15$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst14$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(C),
    .sel(magma_Bit_or_inst1_out),
    .out(Mux2xBit_inst15$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst16$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst15$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(magma_Bit_not_inst0_out),
    .sel(magma_Bits_5_eq_inst18_out),
    .out(Mux2xBit_inst16$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst17$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst16$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(Z),
    .sel(magma_Bits_5_eq_inst19_out),
    .out(Mux2xBit_inst17$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(magma_Bit_or_inst4_out),
    .sel(magma_Bits_5_eq_inst2_out),
    .out(Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(alu),
    .sel(magma_Bits_5_eq_inst3_out),
    .out(Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(magma_Bit_or_inst3_out),
    .sel(magma_Bits_5_eq_inst4_out),
    .out(Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst5$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(magma_Bit_and_inst1_out),
    .sel(magma_Bits_5_eq_inst5_out),
    .out(Mux2xBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst6$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst5$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(magma_Bit_xor_inst1_out),
    .sel(magma_Bits_5_eq_inst6_out),
    .out(Mux2xBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst7$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst6$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(magma_Bit_not_inst6_out),
    .sel(magma_Bits_5_eq_inst7_out),
    .out(Mux2xBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst8$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst7$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(magma_Bit_or_inst2_out),
    .sel(magma_Bits_5_eq_inst8_out),
    .out(Mux2xBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst9$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst8$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(magma_Bit_and_inst0_out),
    .sel(magma_Bits_5_eq_inst9_out),
    .out(Mux2xBit_inst9$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_const #(
    .value(5'h00),
    .width(5)
) const_0_5 (
    .out(const_0_5_out)
);
coreir_const #(
    .value(5'h0a),
    .width(5)
) const_10_5 (
    .out(const_10_5_out)
);
coreir_const #(
    .value(5'h0b),
    .width(5)
) const_11_5 (
    .out(const_11_5_out)
);
coreir_const #(
    .value(5'h0c),
    .width(5)
) const_12_5 (
    .out(const_12_5_out)
);
coreir_const #(
    .value(5'h0d),
    .width(5)
) const_13_5 (
    .out(const_13_5_out)
);
coreir_const #(
    .value(5'h0e),
    .width(5)
) const_14_5 (
    .out(const_14_5_out)
);
coreir_const #(
    .value(5'h0f),
    .width(5)
) const_15_5 (
    .out(const_15_5_out)
);
coreir_const #(
    .value(5'h10),
    .width(5)
) const_16_5 (
    .out(const_16_5_out)
);
coreir_const #(
    .value(5'h11),
    .width(5)
) const_17_5 (
    .out(const_17_5_out)
);
coreir_const #(
    .value(5'h01),
    .width(5)
) const_1_5 (
    .out(const_1_5_out)
);
coreir_const #(
    .value(5'h02),
    .width(5)
) const_2_5 (
    .out(const_2_5_out)
);
coreir_const #(
    .value(5'h03),
    .width(5)
) const_3_5 (
    .out(const_3_5_out)
);
coreir_const #(
    .value(5'h04),
    .width(5)
) const_4_5 (
    .out(const_4_5_out)
);
coreir_const #(
    .value(5'h05),
    .width(5)
) const_5_5 (
    .out(const_5_5_out)
);
coreir_const #(
    .value(5'h06),
    .width(5)
) const_6_5 (
    .out(const_6_5_out)
);
coreir_const #(
    .value(5'h07),
    .width(5)
) const_7_5 (
    .out(const_7_5_out)
);
coreir_const #(
    .value(5'h08),
    .width(5)
) const_8_5 (
    .out(const_8_5_out)
);
coreir_const #(
    .value(5'h09),
    .width(5)
) const_9_5 (
    .out(const_9_5_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(C),
    .in1(magma_Bit_not_inst4_out),
    .out(magma_Bit_and_inst0_out)
);
corebit_and magma_Bit_and_inst1 (
    .in0(magma_Bit_not_inst7_out),
    .in1(magma_Bit_not_inst8_out),
    .out(magma_Bit_and_inst1_out)
);
corebit_and magma_Bit_and_inst2 (
    .in0(magma_Bit_not_inst10_out),
    .in1(magma_Bit_not_inst11_out),
    .out(magma_Bit_and_inst2_out)
);
corebit_and magma_Bit_and_inst3 (
    .in0(N),
    .in1(magma_Bit_not_inst12_out),
    .out(magma_Bit_and_inst3_out)
);
corebit_not magma_Bit_not_inst0 (
    .in(Z),
    .out(magma_Bit_not_inst0_out)
);
corebit_not magma_Bit_not_inst1 (
    .in(C),
    .out(magma_Bit_not_inst1_out)
);
corebit_not magma_Bit_not_inst10 (
    .in(N),
    .out(magma_Bit_not_inst10_out)
);
corebit_not magma_Bit_not_inst11 (
    .in(Z),
    .out(magma_Bit_not_inst11_out)
);
corebit_not magma_Bit_not_inst12 (
    .in(Z),
    .out(magma_Bit_not_inst12_out)
);
corebit_not magma_Bit_not_inst2 (
    .in(N),
    .out(magma_Bit_not_inst2_out)
);
corebit_not magma_Bit_not_inst3 (
    .in(V),
    .out(magma_Bit_not_inst3_out)
);
corebit_not magma_Bit_not_inst4 (
    .in(Z),
    .out(magma_Bit_not_inst4_out)
);
corebit_not magma_Bit_not_inst5 (
    .in(C),
    .out(magma_Bit_not_inst5_out)
);
corebit_not magma_Bit_not_inst6 (
    .in(magma_Bit_xor_inst0_out),
    .out(magma_Bit_not_inst6_out)
);
corebit_not magma_Bit_not_inst7 (
    .in(Z),
    .out(magma_Bit_not_inst7_out)
);
corebit_not magma_Bit_not_inst8 (
    .in(magma_Bit_xor_inst2_out),
    .out(magma_Bit_not_inst8_out)
);
corebit_not magma_Bit_not_inst9 (
    .in(N),
    .out(magma_Bit_not_inst9_out)
);
corebit_or magma_Bit_or_inst0 (
    .in0(magma_Bits_5_eq_inst14_out),
    .in1(magma_Bits_5_eq_inst15_out),
    .out(magma_Bit_or_inst0_out)
);
corebit_or magma_Bit_or_inst1 (
    .in0(magma_Bits_5_eq_inst16_out),
    .in1(magma_Bits_5_eq_inst17_out),
    .out(magma_Bit_or_inst1_out)
);
corebit_or magma_Bit_or_inst2 (
    .in0(magma_Bit_not_inst5_out),
    .in1(Z),
    .out(magma_Bit_or_inst2_out)
);
corebit_or magma_Bit_or_inst3 (
    .in0(Z),
    .in1(magma_Bit_xor_inst3_out),
    .out(magma_Bit_or_inst3_out)
);
corebit_or magma_Bit_or_inst4 (
    .in0(magma_Bit_not_inst9_out),
    .in1(Z),
    .out(magma_Bit_or_inst4_out)
);
corebit_or magma_Bit_or_inst5 (
    .in0(N),
    .in1(Z),
    .out(magma_Bit_or_inst5_out)
);
corebit_xor magma_Bit_xor_inst0 (
    .in0(N),
    .in1(V),
    .out(magma_Bit_xor_inst0_out)
);
corebit_xor magma_Bit_xor_inst1 (
    .in0(N),
    .in1(V),
    .out(magma_Bit_xor_inst1_out)
);
corebit_xor magma_Bit_xor_inst2 (
    .in0(N),
    .in1(V),
    .out(magma_Bit_xor_inst2_out)
);
corebit_xor magma_Bit_xor_inst3 (
    .in0(N),
    .in1(V),
    .out(magma_Bit_xor_inst3_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst0 (
    .in0(code),
    .in1(const_17_5_out),
    .out(magma_Bits_5_eq_inst0_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst1 (
    .in0(code),
    .in1(const_16_5_out),
    .out(magma_Bits_5_eq_inst1_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst10 (
    .in0(code),
    .in1(const_7_5_out),
    .out(magma_Bits_5_eq_inst10_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst11 (
    .in0(code),
    .in1(const_6_5_out),
    .out(magma_Bits_5_eq_inst11_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst12 (
    .in0(code),
    .in1(const_5_5_out),
    .out(magma_Bits_5_eq_inst12_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst13 (
    .in0(code),
    .in1(const_4_5_out),
    .out(magma_Bits_5_eq_inst13_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst14 (
    .in0(code),
    .in1(const_3_5_out),
    .out(magma_Bits_5_eq_inst14_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst15 (
    .in0(code),
    .in1(const_3_5_out),
    .out(magma_Bits_5_eq_inst15_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst16 (
    .in0(code),
    .in1(const_2_5_out),
    .out(magma_Bits_5_eq_inst16_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst17 (
    .in0(code),
    .in1(const_2_5_out),
    .out(magma_Bits_5_eq_inst17_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst18 (
    .in0(code),
    .in1(const_1_5_out),
    .out(magma_Bits_5_eq_inst18_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst19 (
    .in0(code),
    .in1(const_0_5_out),
    .out(magma_Bits_5_eq_inst19_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst2 (
    .in0(code),
    .in1(const_15_5_out),
    .out(magma_Bits_5_eq_inst2_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst3 (
    .in0(code),
    .in1(const_14_5_out),
    .out(magma_Bits_5_eq_inst3_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst4 (
    .in0(code),
    .in1(const_13_5_out),
    .out(magma_Bits_5_eq_inst4_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst5 (
    .in0(code),
    .in1(const_12_5_out),
    .out(magma_Bits_5_eq_inst5_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst6 (
    .in0(code),
    .in1(const_11_5_out),
    .out(magma_Bits_5_eq_inst6_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst7 (
    .in0(code),
    .in1(const_10_5_out),
    .out(magma_Bits_5_eq_inst7_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst8 (
    .in0(code),
    .in1(const_9_5_out),
    .out(magma_Bits_5_eq_inst8_out)
);
coreir_eq #(
    .width(5)
) magma_Bits_5_eq_inst9 (
    .in0(code),
    .in1(const_8_5_out),
    .out(magma_Bits_5_eq_inst9_out)
);
assign O = Mux2xBit_inst17$coreir_commonlib_mux2x1_inst0$_join_out[0];
endmodule

module CB_wen_in_1_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_wen_in_1 (
    input [0:0] I_0,
    input [0:0] I_1,
    input [0:0] I_10,
    input [0:0] I_11,
    input [0:0] I_12,
    input [0:0] I_13,
    input [0:0] I_14,
    input [0:0] I_15,
    input [0:0] I_16,
    input [0:0] I_17,
    input [0:0] I_18,
    input [0:0] I_19,
    input [0:0] I_2,
    input [0:0] I_3,
    input [0:0] I_4,
    input [0:0] I_5,
    input [0:0] I_6,
    input [0:0] I_7,
    input [0:0] I_8,
    input [0:0] I_9,
    output [0:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [4:0] CB_wen_in_1_sel_inst0_O;
wire [0:0] MUX_CB_wen_in_1$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0_out;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [4:0] ZextWrapper_5_32_inst0$self_I_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
CB_wen_in_1_sel CB_wen_in_1_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_wen_in_1_sel_inst0_O)
);
commonlib_muxn__N20__width1 MUX_CB_wen_in_1$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0 (
    .in_data_0(I_0),
    .in_data_1(I_1),
    .in_data_10(I_10),
    .in_data_11(I_11),
    .in_data_12(I_12),
    .in_data_13(I_13),
    .in_data_14(I_14),
    .in_data_15(I_15),
    .in_data_16(I_16),
    .in_data_17(I_17),
    .in_data_18(I_18),
    .in_data_19(I_19),
    .in_data_2(I_2),
    .in_data_3(I_3),
    .in_data_4(I_4),
    .in_data_5(I_5),
    .in_data_6(I_6),
    .in_data_7(I_7),
    .in_data_8(I_8),
    .in_data_9(I_9),
    .in_sel(CB_wen_in_1_sel_inst0_O),
    .out(MUX_CB_wen_in_1$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit5 ZextWrapper_5_32_inst0$self_I (
    .in(config_reg_0_O),
    .out(ZextWrapper_5_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$self_I_out[4:0]};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = MUX_CB_wen_in_1$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0_out;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_wen_in_0_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_wen_in_0 (
    input [0:0] I_0,
    input [0:0] I_1,
    input [0:0] I_10,
    input [0:0] I_11,
    input [0:0] I_12,
    input [0:0] I_13,
    input [0:0] I_14,
    input [0:0] I_15,
    input [0:0] I_16,
    input [0:0] I_17,
    input [0:0] I_18,
    input [0:0] I_19,
    input [0:0] I_2,
    input [0:0] I_3,
    input [0:0] I_4,
    input [0:0] I_5,
    input [0:0] I_6,
    input [0:0] I_7,
    input [0:0] I_8,
    input [0:0] I_9,
    output [0:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [4:0] CB_wen_in_0_sel_inst0_O;
wire [0:0] MUX_CB_wen_in_0$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0_out;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [4:0] ZextWrapper_5_32_inst0$self_I_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
CB_wen_in_0_sel CB_wen_in_0_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_wen_in_0_sel_inst0_O)
);
commonlib_muxn__N20__width1 MUX_CB_wen_in_0$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0 (
    .in_data_0(I_0),
    .in_data_1(I_1),
    .in_data_10(I_10),
    .in_data_11(I_11),
    .in_data_12(I_12),
    .in_data_13(I_13),
    .in_data_14(I_14),
    .in_data_15(I_15),
    .in_data_16(I_16),
    .in_data_17(I_17),
    .in_data_18(I_18),
    .in_data_19(I_19),
    .in_data_2(I_2),
    .in_data_3(I_3),
    .in_data_4(I_4),
    .in_data_5(I_5),
    .in_data_6(I_6),
    .in_data_7(I_7),
    .in_data_8(I_8),
    .in_data_9(I_9),
    .in_sel(CB_wen_in_0_sel_inst0_O),
    .out(MUX_CB_wen_in_0$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit5 ZextWrapper_5_32_inst0$self_I (
    .in(config_reg_0_O),
    .out(ZextWrapper_5_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$self_I_out[4:0]};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = MUX_CB_wen_in_0$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0_out;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_ren_in_1_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_ren_in_1 (
    input [0:0] I_0,
    input [0:0] I_1,
    input [0:0] I_10,
    input [0:0] I_11,
    input [0:0] I_12,
    input [0:0] I_13,
    input [0:0] I_14,
    input [0:0] I_15,
    input [0:0] I_16,
    input [0:0] I_17,
    input [0:0] I_18,
    input [0:0] I_19,
    input [0:0] I_2,
    input [0:0] I_3,
    input [0:0] I_4,
    input [0:0] I_5,
    input [0:0] I_6,
    input [0:0] I_7,
    input [0:0] I_8,
    input [0:0] I_9,
    output [0:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [4:0] CB_ren_in_1_sel_inst0_O;
wire [0:0] MUX_CB_ren_in_1$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0_out;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [4:0] ZextWrapper_5_32_inst0$self_I_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
CB_ren_in_1_sel CB_ren_in_1_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_ren_in_1_sel_inst0_O)
);
commonlib_muxn__N20__width1 MUX_CB_ren_in_1$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0 (
    .in_data_0(I_0),
    .in_data_1(I_1),
    .in_data_10(I_10),
    .in_data_11(I_11),
    .in_data_12(I_12),
    .in_data_13(I_13),
    .in_data_14(I_14),
    .in_data_15(I_15),
    .in_data_16(I_16),
    .in_data_17(I_17),
    .in_data_18(I_18),
    .in_data_19(I_19),
    .in_data_2(I_2),
    .in_data_3(I_3),
    .in_data_4(I_4),
    .in_data_5(I_5),
    .in_data_6(I_6),
    .in_data_7(I_7),
    .in_data_8(I_8),
    .in_data_9(I_9),
    .in_sel(CB_ren_in_1_sel_inst0_O),
    .out(MUX_CB_ren_in_1$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit5 ZextWrapper_5_32_inst0$self_I (
    .in(config_reg_0_O),
    .out(ZextWrapper_5_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$self_I_out[4:0]};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = MUX_CB_ren_in_1$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0_out;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_ren_in_0_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_ren_in_0 (
    input [0:0] I_0,
    input [0:0] I_1,
    input [0:0] I_10,
    input [0:0] I_11,
    input [0:0] I_12,
    input [0:0] I_13,
    input [0:0] I_14,
    input [0:0] I_15,
    input [0:0] I_16,
    input [0:0] I_17,
    input [0:0] I_18,
    input [0:0] I_19,
    input [0:0] I_2,
    input [0:0] I_3,
    input [0:0] I_4,
    input [0:0] I_5,
    input [0:0] I_6,
    input [0:0] I_7,
    input [0:0] I_8,
    input [0:0] I_9,
    output [0:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [4:0] CB_ren_in_0_sel_inst0_O;
wire [0:0] MUX_CB_ren_in_0$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0_out;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [4:0] ZextWrapper_5_32_inst0$self_I_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
CB_ren_in_0_sel CB_ren_in_0_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_ren_in_0_sel_inst0_O)
);
commonlib_muxn__N20__width1 MUX_CB_ren_in_0$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0 (
    .in_data_0(I_0),
    .in_data_1(I_1),
    .in_data_10(I_10),
    .in_data_11(I_11),
    .in_data_12(I_12),
    .in_data_13(I_13),
    .in_data_14(I_14),
    .in_data_15(I_15),
    .in_data_16(I_16),
    .in_data_17(I_17),
    .in_data_18(I_18),
    .in_data_19(I_19),
    .in_data_2(I_2),
    .in_data_3(I_3),
    .in_data_4(I_4),
    .in_data_5(I_5),
    .in_data_6(I_6),
    .in_data_7(I_7),
    .in_data_8(I_8),
    .in_data_9(I_9),
    .in_sel(CB_ren_in_0_sel_inst0_O),
    .out(MUX_CB_ren_in_0$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit5 ZextWrapper_5_32_inst0$self_I (
    .in(config_reg_0_O),
    .out(ZextWrapper_5_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$self_I_out[4:0]};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = MUX_CB_ren_in_0$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0_out;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_inputs5_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_inputs5 (
    input [0:0] I_0,
    input [0:0] I_1,
    input [0:0] I_10,
    input [0:0] I_11,
    input [0:0] I_12,
    input [0:0] I_13,
    input [0:0] I_14,
    input [0:0] I_15,
    input [0:0] I_16,
    input [0:0] I_17,
    input [0:0] I_18,
    input [0:0] I_19,
    input [0:0] I_2,
    input [0:0] I_3,
    input [0:0] I_4,
    input [0:0] I_5,
    input [0:0] I_6,
    input [0:0] I_7,
    input [0:0] I_8,
    input [0:0] I_9,
    output [0:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [4:0] CB_inputs5_sel_inst0_O;
wire [0:0] MUX_CB_inputs5$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0_out;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [4:0] ZextWrapper_5_32_inst0$self_I_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
CB_inputs5_sel CB_inputs5_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_inputs5_sel_inst0_O)
);
commonlib_muxn__N20__width1 MUX_CB_inputs5$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0 (
    .in_data_0(I_0),
    .in_data_1(I_1),
    .in_data_10(I_10),
    .in_data_11(I_11),
    .in_data_12(I_12),
    .in_data_13(I_13),
    .in_data_14(I_14),
    .in_data_15(I_15),
    .in_data_16(I_16),
    .in_data_17(I_17),
    .in_data_18(I_18),
    .in_data_19(I_19),
    .in_data_2(I_2),
    .in_data_3(I_3),
    .in_data_4(I_4),
    .in_data_5(I_5),
    .in_data_6(I_6),
    .in_data_7(I_7),
    .in_data_8(I_8),
    .in_data_9(I_9),
    .in_sel(CB_inputs5_sel_inst0_O),
    .out(MUX_CB_inputs5$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit5 ZextWrapper_5_32_inst0$self_I (
    .in(config_reg_0_O),
    .out(ZextWrapper_5_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$self_I_out[4:0]};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = MUX_CB_inputs5$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0_out;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_inputs4_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_inputs4 (
    input [0:0] I_0,
    input [0:0] I_1,
    input [0:0] I_10,
    input [0:0] I_11,
    input [0:0] I_12,
    input [0:0] I_13,
    input [0:0] I_14,
    input [0:0] I_15,
    input [0:0] I_16,
    input [0:0] I_17,
    input [0:0] I_18,
    input [0:0] I_19,
    input [0:0] I_2,
    input [0:0] I_3,
    input [0:0] I_4,
    input [0:0] I_5,
    input [0:0] I_6,
    input [0:0] I_7,
    input [0:0] I_8,
    input [0:0] I_9,
    output [0:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [4:0] CB_inputs4_sel_inst0_O;
wire [0:0] MUX_CB_inputs4$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0_out;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [4:0] ZextWrapper_5_32_inst0$self_I_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
CB_inputs4_sel CB_inputs4_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_inputs4_sel_inst0_O)
);
commonlib_muxn__N20__width1 MUX_CB_inputs4$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0 (
    .in_data_0(I_0),
    .in_data_1(I_1),
    .in_data_10(I_10),
    .in_data_11(I_11),
    .in_data_12(I_12),
    .in_data_13(I_13),
    .in_data_14(I_14),
    .in_data_15(I_15),
    .in_data_16(I_16),
    .in_data_17(I_17),
    .in_data_18(I_18),
    .in_data_19(I_19),
    .in_data_2(I_2),
    .in_data_3(I_3),
    .in_data_4(I_4),
    .in_data_5(I_5),
    .in_data_6(I_6),
    .in_data_7(I_7),
    .in_data_8(I_8),
    .in_data_9(I_9),
    .in_sel(CB_inputs4_sel_inst0_O),
    .out(MUX_CB_inputs4$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit5 ZextWrapper_5_32_inst0$self_I (
    .in(config_reg_0_O),
    .out(ZextWrapper_5_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$self_I_out[4:0]};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = MUX_CB_inputs4$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0_out;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_inputs3_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_inputs3 (
    input [0:0] I_0,
    input [0:0] I_1,
    input [0:0] I_10,
    input [0:0] I_11,
    input [0:0] I_12,
    input [0:0] I_13,
    input [0:0] I_14,
    input [0:0] I_15,
    input [0:0] I_16,
    input [0:0] I_17,
    input [0:0] I_18,
    input [0:0] I_19,
    input [0:0] I_2,
    input [0:0] I_3,
    input [0:0] I_4,
    input [0:0] I_5,
    input [0:0] I_6,
    input [0:0] I_7,
    input [0:0] I_8,
    input [0:0] I_9,
    output [0:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [4:0] CB_inputs3_sel_inst0_O;
wire [0:0] MUX_CB_inputs3$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0_out;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [4:0] ZextWrapper_5_32_inst0$self_I_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
CB_inputs3_sel CB_inputs3_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_inputs3_sel_inst0_O)
);
commonlib_muxn__N20__width1 MUX_CB_inputs3$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0 (
    .in_data_0(I_0),
    .in_data_1(I_1),
    .in_data_10(I_10),
    .in_data_11(I_11),
    .in_data_12(I_12),
    .in_data_13(I_13),
    .in_data_14(I_14),
    .in_data_15(I_15),
    .in_data_16(I_16),
    .in_data_17(I_17),
    .in_data_18(I_18),
    .in_data_19(I_19),
    .in_data_2(I_2),
    .in_data_3(I_3),
    .in_data_4(I_4),
    .in_data_5(I_5),
    .in_data_6(I_6),
    .in_data_7(I_7),
    .in_data_8(I_8),
    .in_data_9(I_9),
    .in_sel(CB_inputs3_sel_inst0_O),
    .out(MUX_CB_inputs3$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit5 ZextWrapper_5_32_inst0$self_I (
    .in(config_reg_0_O),
    .out(ZextWrapper_5_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$self_I_out[4:0]};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = MUX_CB_inputs3$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0_out;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_inputs2_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_inputs2 (
    input [15:0] I_0,
    input [15:0] I_1,
    input [15:0] I_10,
    input [15:0] I_11,
    input [15:0] I_12,
    input [15:0] I_13,
    input [15:0] I_14,
    input [15:0] I_15,
    input [15:0] I_16,
    input [15:0] I_17,
    input [15:0] I_18,
    input [15:0] I_19,
    input [15:0] I_2,
    input [15:0] I_3,
    input [15:0] I_4,
    input [15:0] I_5,
    input [15:0] I_6,
    input [15:0] I_7,
    input [15:0] I_8,
    input [15:0] I_9,
    output [15:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [4:0] CB_inputs2_sel_inst0_O;
wire [15:0] MUX_CB_inputs2$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [4:0] ZextWrapper_5_32_inst0$self_I_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
CB_inputs2_sel CB_inputs2_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_inputs2_sel_inst0_O)
);
commonlib_muxn__N20__width16 MUX_CB_inputs2$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0 (
    .in_data_0(I_0),
    .in_data_1(I_1),
    .in_data_10(I_10),
    .in_data_11(I_11),
    .in_data_12(I_12),
    .in_data_13(I_13),
    .in_data_14(I_14),
    .in_data_15(I_15),
    .in_data_16(I_16),
    .in_data_17(I_17),
    .in_data_18(I_18),
    .in_data_19(I_19),
    .in_data_2(I_2),
    .in_data_3(I_3),
    .in_data_4(I_4),
    .in_data_5(I_5),
    .in_data_6(I_6),
    .in_data_7(I_7),
    .in_data_8(I_8),
    .in_data_9(I_9),
    .in_sel(CB_inputs2_sel_inst0_O),
    .out(MUX_CB_inputs2$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit5 ZextWrapper_5_32_inst0$self_I (
    .in(config_reg_0_O),
    .out(ZextWrapper_5_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$self_I_out[4:0]};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = MUX_CB_inputs2$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_inputs1_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_inputs1 (
    input [15:0] I_0,
    input [15:0] I_1,
    input [15:0] I_10,
    input [15:0] I_11,
    input [15:0] I_12,
    input [15:0] I_13,
    input [15:0] I_14,
    input [15:0] I_15,
    input [15:0] I_16,
    input [15:0] I_17,
    input [15:0] I_18,
    input [15:0] I_19,
    input [15:0] I_2,
    input [15:0] I_3,
    input [15:0] I_4,
    input [15:0] I_5,
    input [15:0] I_6,
    input [15:0] I_7,
    input [15:0] I_8,
    input [15:0] I_9,
    output [15:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [4:0] CB_inputs1_sel_inst0_O;
wire [15:0] MUX_CB_inputs1$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [4:0] ZextWrapper_5_32_inst0$self_I_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
CB_inputs1_sel CB_inputs1_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_inputs1_sel_inst0_O)
);
commonlib_muxn__N20__width16 MUX_CB_inputs1$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0 (
    .in_data_0(I_0),
    .in_data_1(I_1),
    .in_data_10(I_10),
    .in_data_11(I_11),
    .in_data_12(I_12),
    .in_data_13(I_13),
    .in_data_14(I_14),
    .in_data_15(I_15),
    .in_data_16(I_16),
    .in_data_17(I_17),
    .in_data_18(I_18),
    .in_data_19(I_19),
    .in_data_2(I_2),
    .in_data_3(I_3),
    .in_data_4(I_4),
    .in_data_5(I_5),
    .in_data_6(I_6),
    .in_data_7(I_7),
    .in_data_8(I_8),
    .in_data_9(I_9),
    .in_sel(CB_inputs1_sel_inst0_O),
    .out(MUX_CB_inputs1$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit5 ZextWrapper_5_32_inst0$self_I (
    .in(config_reg_0_O),
    .out(ZextWrapper_5_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$self_I_out[4:0]};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = MUX_CB_inputs1$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_inputs0_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_inputs0 (
    input [15:0] I_0,
    input [15:0] I_1,
    input [15:0] I_10,
    input [15:0] I_11,
    input [15:0] I_12,
    input [15:0] I_13,
    input [15:0] I_14,
    input [15:0] I_15,
    input [15:0] I_16,
    input [15:0] I_17,
    input [15:0] I_18,
    input [15:0] I_19,
    input [15:0] I_2,
    input [15:0] I_3,
    input [15:0] I_4,
    input [15:0] I_5,
    input [15:0] I_6,
    input [15:0] I_7,
    input [15:0] I_8,
    input [15:0] I_9,
    output [15:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [4:0] CB_inputs0_sel_inst0_O;
wire [15:0] MUX_CB_inputs0$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [4:0] ZextWrapper_5_32_inst0$self_I_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
CB_inputs0_sel CB_inputs0_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_inputs0_sel_inst0_O)
);
commonlib_muxn__N20__width16 MUX_CB_inputs0$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0 (
    .in_data_0(I_0),
    .in_data_1(I_1),
    .in_data_10(I_10),
    .in_data_11(I_11),
    .in_data_12(I_12),
    .in_data_13(I_13),
    .in_data_14(I_14),
    .in_data_15(I_15),
    .in_data_16(I_16),
    .in_data_17(I_17),
    .in_data_18(I_18),
    .in_data_19(I_19),
    .in_data_2(I_2),
    .in_data_3(I_3),
    .in_data_4(I_4),
    .in_data_5(I_5),
    .in_data_6(I_6),
    .in_data_7(I_7),
    .in_data_8(I_8),
    .in_data_9(I_9),
    .in_sel(CB_inputs0_sel_inst0_O),
    .out(MUX_CB_inputs0$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit5 ZextWrapper_5_32_inst0$self_I (
    .in(config_reg_0_O),
    .out(ZextWrapper_5_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$self_I_out[4:0]};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = MUX_CB_inputs0$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_flush_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_flush (
    input [0:0] I_0,
    input [0:0] I_1,
    input [0:0] I_10,
    input [0:0] I_11,
    input [0:0] I_12,
    input [0:0] I_13,
    input [0:0] I_14,
    input [0:0] I_15,
    input [0:0] I_16,
    input [0:0] I_17,
    input [0:0] I_18,
    input [0:0] I_19,
    input [0:0] I_2,
    input [0:0] I_3,
    input [0:0] I_4,
    input [0:0] I_5,
    input [0:0] I_6,
    input [0:0] I_7,
    input [0:0] I_8,
    input [0:0] I_9,
    output [0:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [4:0] CB_flush_sel_inst0_O;
wire [0:0] MUX_CB_flush$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0_out;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [4:0] ZextWrapper_5_32_inst0$self_I_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
CB_flush_sel CB_flush_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_flush_sel_inst0_O)
);
commonlib_muxn__N20__width1 MUX_CB_flush$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0 (
    .in_data_0(I_0),
    .in_data_1(I_1),
    .in_data_10(I_10),
    .in_data_11(I_11),
    .in_data_12(I_12),
    .in_data_13(I_13),
    .in_data_14(I_14),
    .in_data_15(I_15),
    .in_data_16(I_16),
    .in_data_17(I_17),
    .in_data_18(I_18),
    .in_data_19(I_19),
    .in_data_2(I_2),
    .in_data_3(I_3),
    .in_data_4(I_4),
    .in_data_5(I_5),
    .in_data_6(I_6),
    .in_data_7(I_7),
    .in_data_8(I_8),
    .in_data_9(I_9),
    .in_sel(CB_flush_sel_inst0_O),
    .out(MUX_CB_flush$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit5 ZextWrapper_5_32_inst0$self_I (
    .in(config_reg_0_O),
    .out(ZextWrapper_5_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$self_I_out[4:0]};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = MUX_CB_flush$Mux20x1_inst0$coreir_commonlib_mux20x1_inst0_out;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_data_in_1_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_data_in_1 (
    input [15:0] I_0,
    input [15:0] I_1,
    input [15:0] I_10,
    input [15:0] I_11,
    input [15:0] I_12,
    input [15:0] I_13,
    input [15:0] I_14,
    input [15:0] I_15,
    input [15:0] I_16,
    input [15:0] I_17,
    input [15:0] I_18,
    input [15:0] I_19,
    input [15:0] I_2,
    input [15:0] I_3,
    input [15:0] I_4,
    input [15:0] I_5,
    input [15:0] I_6,
    input [15:0] I_7,
    input [15:0] I_8,
    input [15:0] I_9,
    output [15:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [4:0] CB_data_in_1_sel_inst0_O;
wire [15:0] MUX_CB_data_in_1$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [4:0] ZextWrapper_5_32_inst0$self_I_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
CB_data_in_1_sel CB_data_in_1_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_data_in_1_sel_inst0_O)
);
commonlib_muxn__N20__width16 MUX_CB_data_in_1$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0 (
    .in_data_0(I_0),
    .in_data_1(I_1),
    .in_data_10(I_10),
    .in_data_11(I_11),
    .in_data_12(I_12),
    .in_data_13(I_13),
    .in_data_14(I_14),
    .in_data_15(I_15),
    .in_data_16(I_16),
    .in_data_17(I_17),
    .in_data_18(I_18),
    .in_data_19(I_19),
    .in_data_2(I_2),
    .in_data_3(I_3),
    .in_data_4(I_4),
    .in_data_5(I_5),
    .in_data_6(I_6),
    .in_data_7(I_7),
    .in_data_8(I_8),
    .in_data_9(I_9),
    .in_sel(CB_data_in_1_sel_inst0_O),
    .out(MUX_CB_data_in_1$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit5 ZextWrapper_5_32_inst0$self_I (
    .in(config_reg_0_O),
    .out(ZextWrapper_5_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$self_I_out[4:0]};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = MUX_CB_data_in_1$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_data_in_0_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_data_in_0 (
    input [15:0] I_0,
    input [15:0] I_1,
    input [15:0] I_10,
    input [15:0] I_11,
    input [15:0] I_12,
    input [15:0] I_13,
    input [15:0] I_14,
    input [15:0] I_15,
    input [15:0] I_16,
    input [15:0] I_17,
    input [15:0] I_18,
    input [15:0] I_19,
    input [15:0] I_2,
    input [15:0] I_3,
    input [15:0] I_4,
    input [15:0] I_5,
    input [15:0] I_6,
    input [15:0] I_7,
    input [15:0] I_8,
    input [15:0] I_9,
    output [15:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [4:0] CB_data_in_0_sel_inst0_O;
wire [15:0] MUX_CB_data_in_0$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [4:0] ZextWrapper_5_32_inst0$self_I_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
CB_data_in_0_sel CB_data_in_0_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_data_in_0_sel_inst0_O)
);
commonlib_muxn__N20__width16 MUX_CB_data_in_0$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0 (
    .in_data_0(I_0),
    .in_data_1(I_1),
    .in_data_10(I_10),
    .in_data_11(I_11),
    .in_data_12(I_12),
    .in_data_13(I_13),
    .in_data_14(I_14),
    .in_data_15(I_15),
    .in_data_16(I_16),
    .in_data_17(I_17),
    .in_data_18(I_18),
    .in_data_19(I_19),
    .in_data_2(I_2),
    .in_data_3(I_3),
    .in_data_4(I_4),
    .in_data_5(I_5),
    .in_data_6(I_6),
    .in_data_7(I_7),
    .in_data_8(I_8),
    .in_data_9(I_9),
    .in_sel(CB_data_in_0_sel_inst0_O),
    .out(MUX_CB_data_in_0$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit5 ZextWrapper_5_32_inst0$self_I (
    .in(config_reg_0_O),
    .out(ZextWrapper_5_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$self_I_out[4:0]};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = MUX_CB_data_in_0$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_chain_data_in_1_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_chain_data_in_1 (
    input [15:0] I_0,
    input [15:0] I_1,
    input [15:0] I_10,
    input [15:0] I_11,
    input [15:0] I_12,
    input [15:0] I_13,
    input [15:0] I_14,
    input [15:0] I_15,
    input [15:0] I_16,
    input [15:0] I_17,
    input [15:0] I_18,
    input [15:0] I_19,
    input [15:0] I_2,
    input [15:0] I_3,
    input [15:0] I_4,
    input [15:0] I_5,
    input [15:0] I_6,
    input [15:0] I_7,
    input [15:0] I_8,
    input [15:0] I_9,
    output [15:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [4:0] CB_chain_data_in_1_sel_inst0_O;
wire [15:0] MUX_CB_chain_data_in_1$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [4:0] ZextWrapper_5_32_inst0$self_I_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
CB_chain_data_in_1_sel CB_chain_data_in_1_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_chain_data_in_1_sel_inst0_O)
);
commonlib_muxn__N20__width16 MUX_CB_chain_data_in_1$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0 (
    .in_data_0(I_0),
    .in_data_1(I_1),
    .in_data_10(I_10),
    .in_data_11(I_11),
    .in_data_12(I_12),
    .in_data_13(I_13),
    .in_data_14(I_14),
    .in_data_15(I_15),
    .in_data_16(I_16),
    .in_data_17(I_17),
    .in_data_18(I_18),
    .in_data_19(I_19),
    .in_data_2(I_2),
    .in_data_3(I_3),
    .in_data_4(I_4),
    .in_data_5(I_5),
    .in_data_6(I_6),
    .in_data_7(I_7),
    .in_data_8(I_8),
    .in_data_9(I_9),
    .in_sel(CB_chain_data_in_1_sel_inst0_O),
    .out(MUX_CB_chain_data_in_1$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit5 ZextWrapper_5_32_inst0$self_I (
    .in(config_reg_0_O),
    .out(ZextWrapper_5_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$self_I_out[4:0]};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = MUX_CB_chain_data_in_1$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_chain_data_in_0_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_chain_data_in_0 (
    input [15:0] I_0,
    input [15:0] I_1,
    input [15:0] I_10,
    input [15:0] I_11,
    input [15:0] I_12,
    input [15:0] I_13,
    input [15:0] I_14,
    input [15:0] I_15,
    input [15:0] I_16,
    input [15:0] I_17,
    input [15:0] I_18,
    input [15:0] I_19,
    input [15:0] I_2,
    input [15:0] I_3,
    input [15:0] I_4,
    input [15:0] I_5,
    input [15:0] I_6,
    input [15:0] I_7,
    input [15:0] I_8,
    input [15:0] I_9,
    output [15:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [4:0] CB_chain_data_in_0_sel_inst0_O;
wire [15:0] MUX_CB_chain_data_in_0$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [4:0] ZextWrapper_5_32_inst0$self_I_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
CB_chain_data_in_0_sel CB_chain_data_in_0_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_chain_data_in_0_sel_inst0_O)
);
commonlib_muxn__N20__width16 MUX_CB_chain_data_in_0$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0 (
    .in_data_0(I_0),
    .in_data_1(I_1),
    .in_data_10(I_10),
    .in_data_11(I_11),
    .in_data_12(I_12),
    .in_data_13(I_13),
    .in_data_14(I_14),
    .in_data_15(I_15),
    .in_data_16(I_16),
    .in_data_17(I_17),
    .in_data_18(I_18),
    .in_data_19(I_19),
    .in_data_2(I_2),
    .in_data_3(I_3),
    .in_data_4(I_4),
    .in_data_5(I_5),
    .in_data_6(I_6),
    .in_data_7(I_7),
    .in_data_8(I_8),
    .in_data_9(I_9),
    .in_sel(CB_chain_data_in_0_sel_inst0_O),
    .out(MUX_CB_chain_data_in_0$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit5 ZextWrapper_5_32_inst0$self_I (
    .in(config_reg_0_O),
    .out(ZextWrapper_5_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$self_I_out[4:0]};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = MUX_CB_chain_data_in_0$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_addr_in_1_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_addr_in_1 (
    input [15:0] I_0,
    input [15:0] I_1,
    input [15:0] I_10,
    input [15:0] I_11,
    input [15:0] I_12,
    input [15:0] I_13,
    input [15:0] I_14,
    input [15:0] I_15,
    input [15:0] I_16,
    input [15:0] I_17,
    input [15:0] I_18,
    input [15:0] I_19,
    input [15:0] I_2,
    input [15:0] I_3,
    input [15:0] I_4,
    input [15:0] I_5,
    input [15:0] I_6,
    input [15:0] I_7,
    input [15:0] I_8,
    input [15:0] I_9,
    output [15:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [4:0] CB_addr_in_1_sel_inst0_O;
wire [15:0] MUX_CB_addr_in_1$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [4:0] ZextWrapper_5_32_inst0$self_I_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
CB_addr_in_1_sel CB_addr_in_1_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_addr_in_1_sel_inst0_O)
);
commonlib_muxn__N20__width16 MUX_CB_addr_in_1$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0 (
    .in_data_0(I_0),
    .in_data_1(I_1),
    .in_data_10(I_10),
    .in_data_11(I_11),
    .in_data_12(I_12),
    .in_data_13(I_13),
    .in_data_14(I_14),
    .in_data_15(I_15),
    .in_data_16(I_16),
    .in_data_17(I_17),
    .in_data_18(I_18),
    .in_data_19(I_19),
    .in_data_2(I_2),
    .in_data_3(I_3),
    .in_data_4(I_4),
    .in_data_5(I_5),
    .in_data_6(I_6),
    .in_data_7(I_7),
    .in_data_8(I_8),
    .in_data_9(I_9),
    .in_sel(CB_addr_in_1_sel_inst0_O),
    .out(MUX_CB_addr_in_1$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit5 ZextWrapper_5_32_inst0$self_I (
    .in(config_reg_0_O),
    .out(ZextWrapper_5_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$self_I_out[4:0]};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = MUX_CB_addr_in_1$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module CB_addr_in_0_sel (
    input [4:0] I,
    output [4:0] O
);
assign O = I;
endmodule

module CB_addr_in_0 (
    input [15:0] I_0,
    input [15:0] I_1,
    input [15:0] I_10,
    input [15:0] I_11,
    input [15:0] I_12,
    input [15:0] I_13,
    input [15:0] I_14,
    input [15:0] I_15,
    input [15:0] I_16,
    input [15:0] I_17,
    input [15:0] I_18,
    input [15:0] I_19,
    input [15:0] I_2,
    input [15:0] I_3,
    input [15:0] I_4,
    input [15:0] I_5,
    input [15:0] I_6,
    input [15:0] I_7,
    input [15:0] I_8,
    input [15:0] I_9,
    output [15:0] O,
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    output [31:0] read_config_data,
    input reset
);
wire [4:0] CB_addr_in_0_sel_inst0_O;
wire [15:0] MUX_CB_addr_in_0$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out;
wire ZextWrapper_5_32_inst0$bit_const_0_None_out;
wire [4:0] ZextWrapper_5_32_inst0$self_I_out;
wire [31:0] ZextWrapper_5_32_inst0$self_O_in;
wire [4:0] config_reg_0_O;
CB_addr_in_0_sel CB_addr_in_0_sel_inst0 (
    .I(config_reg_0_O),
    .O(CB_addr_in_0_sel_inst0_O)
);
commonlib_muxn__N20__width16 MUX_CB_addr_in_0$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0 (
    .in_data_0(I_0),
    .in_data_1(I_1),
    .in_data_10(I_10),
    .in_data_11(I_11),
    .in_data_12(I_12),
    .in_data_13(I_13),
    .in_data_14(I_14),
    .in_data_15(I_15),
    .in_data_16(I_16),
    .in_data_17(I_17),
    .in_data_18(I_18),
    .in_data_19(I_19),
    .in_data_2(I_2),
    .in_data_3(I_3),
    .in_data_4(I_4),
    .in_data_5(I_5),
    .in_data_6(I_6),
    .in_data_7(I_7),
    .in_data_8(I_8),
    .in_data_9(I_9),
    .in_sel(CB_addr_in_0_sel_inst0_O),
    .out(MUX_CB_addr_in_0$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out)
);
corebit_const #(
    .value(1'b0)
) ZextWrapper_5_32_inst0$bit_const_0_None (
    .out(ZextWrapper_5_32_inst0$bit_const_0_None_out)
);
mantle_wire__typeBit5 ZextWrapper_5_32_inst0$self_I (
    .in(config_reg_0_O),
    .out(ZextWrapper_5_32_inst0$self_I_out)
);
wire [31:0] ZextWrapper_5_32_inst0$self_O_out;
assign ZextWrapper_5_32_inst0$self_O_out = {ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$bit_const_0_None_out,ZextWrapper_5_32_inst0$self_I_out[4:0]};
mantle_wire__typeBitIn32 ZextWrapper_5_32_inst0$self_O (
    .in(ZextWrapper_5_32_inst0$self_O_in),
    .out(ZextWrapper_5_32_inst0$self_O_out)
);
ConfigRegister_5_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
assign O = MUX_CB_addr_in_0$Mux20x16_inst0$coreir_commonlib_mux20x16_inst0_out;
assign read_config_data = ZextWrapper_5_32_inst0$self_O_in;
endmodule

module Tile_MemCore (
    input [0:0] SB_T0_EAST_SB_IN_B1,
    input [15:0] SB_T0_EAST_SB_IN_B16,
    output [0:0] SB_T0_EAST_SB_OUT_B1,
    output [15:0] SB_T0_EAST_SB_OUT_B16,
    input [0:0] SB_T0_NORTH_SB_IN_B1,
    input [15:0] SB_T0_NORTH_SB_IN_B16,
    output [0:0] SB_T0_NORTH_SB_OUT_B1,
    output [15:0] SB_T0_NORTH_SB_OUT_B16,
    input [0:0] SB_T0_SOUTH_SB_IN_B1,
    input [15:0] SB_T0_SOUTH_SB_IN_B16,
    output [0:0] SB_T0_SOUTH_SB_OUT_B1,
    output [15:0] SB_T0_SOUTH_SB_OUT_B16,
    input [0:0] SB_T0_WEST_SB_IN_B1,
    input [15:0] SB_T0_WEST_SB_IN_B16,
    output [0:0] SB_T0_WEST_SB_OUT_B1,
    output [15:0] SB_T0_WEST_SB_OUT_B16,
    input [0:0] SB_T1_EAST_SB_IN_B1,
    input [15:0] SB_T1_EAST_SB_IN_B16,
    output [0:0] SB_T1_EAST_SB_OUT_B1,
    output [15:0] SB_T1_EAST_SB_OUT_B16,
    input [0:0] SB_T1_NORTH_SB_IN_B1,
    input [15:0] SB_T1_NORTH_SB_IN_B16,
    output [0:0] SB_T1_NORTH_SB_OUT_B1,
    output [15:0] SB_T1_NORTH_SB_OUT_B16,
    input [0:0] SB_T1_SOUTH_SB_IN_B1,
    input [15:0] SB_T1_SOUTH_SB_IN_B16,
    output [0:0] SB_T1_SOUTH_SB_OUT_B1,
    output [15:0] SB_T1_SOUTH_SB_OUT_B16,
    input [0:0] SB_T1_WEST_SB_IN_B1,
    input [15:0] SB_T1_WEST_SB_IN_B16,
    output [0:0] SB_T1_WEST_SB_OUT_B1,
    output [15:0] SB_T1_WEST_SB_OUT_B16,
    input [0:0] SB_T2_EAST_SB_IN_B1,
    input [15:0] SB_T2_EAST_SB_IN_B16,
    output [0:0] SB_T2_EAST_SB_OUT_B1,
    output [15:0] SB_T2_EAST_SB_OUT_B16,
    input [0:0] SB_T2_NORTH_SB_IN_B1,
    input [15:0] SB_T2_NORTH_SB_IN_B16,
    output [0:0] SB_T2_NORTH_SB_OUT_B1,
    output [15:0] SB_T2_NORTH_SB_OUT_B16,
    input [0:0] SB_T2_SOUTH_SB_IN_B1,
    input [15:0] SB_T2_SOUTH_SB_IN_B16,
    output [0:0] SB_T2_SOUTH_SB_OUT_B1,
    output [15:0] SB_T2_SOUTH_SB_OUT_B16,
    input [0:0] SB_T2_WEST_SB_IN_B1,
    input [15:0] SB_T2_WEST_SB_IN_B16,
    output [0:0] SB_T2_WEST_SB_OUT_B1,
    output [15:0] SB_T2_WEST_SB_OUT_B16,
    input [0:0] SB_T3_EAST_SB_IN_B1,
    input [15:0] SB_T3_EAST_SB_IN_B16,
    output [0:0] SB_T3_EAST_SB_OUT_B1,
    output [15:0] SB_T3_EAST_SB_OUT_B16,
    input [0:0] SB_T3_NORTH_SB_IN_B1,
    input [15:0] SB_T3_NORTH_SB_IN_B16,
    output [0:0] SB_T3_NORTH_SB_OUT_B1,
    output [15:0] SB_T3_NORTH_SB_OUT_B16,
    input [0:0] SB_T3_SOUTH_SB_IN_B1,
    input [15:0] SB_T3_SOUTH_SB_IN_B16,
    output [0:0] SB_T3_SOUTH_SB_OUT_B1,
    output [15:0] SB_T3_SOUTH_SB_OUT_B16,
    input [0:0] SB_T3_WEST_SB_IN_B1,
    input [15:0] SB_T3_WEST_SB_IN_B16,
    output [0:0] SB_T3_WEST_SB_OUT_B1,
    output [15:0] SB_T3_WEST_SB_OUT_B16,
    input [0:0] SB_T4_EAST_SB_IN_B1,
    input [15:0] SB_T4_EAST_SB_IN_B16,
    output [0:0] SB_T4_EAST_SB_OUT_B1,
    output [15:0] SB_T4_EAST_SB_OUT_B16,
    input [0:0] SB_T4_NORTH_SB_IN_B1,
    input [15:0] SB_T4_NORTH_SB_IN_B16,
    output [0:0] SB_T4_NORTH_SB_OUT_B1,
    output [15:0] SB_T4_NORTH_SB_OUT_B16,
    input [0:0] SB_T4_SOUTH_SB_IN_B1,
    input [15:0] SB_T4_SOUTH_SB_IN_B16,
    output [0:0] SB_T4_SOUTH_SB_OUT_B1,
    output [15:0] SB_T4_SOUTH_SB_OUT_B16,
    input [0:0] SB_T4_WEST_SB_IN_B1,
    input [15:0] SB_T4_WEST_SB_IN_B16,
    output [0:0] SB_T4_WEST_SB_OUT_B1,
    output [15:0] SB_T4_WEST_SB_OUT_B16,
    input clk,
    output clk_out,
    input [31:0] config_config_addr,
    input [31:0] config_config_data,
    output [31:0] config_out_config_addr,
    output [31:0] config_out_config_data,
    output [0:0] config_out_read,
    output [0:0] config_out_write,
    input [0:0] config_read,
    input [0:0] config_write,
    output [8:0] hi,
    output [7:0] lo,
    output [31:0] read_config_data,
    input [31:0] read_config_data_in,
    input reset,
    output reset_out,
    input [0:0] stall,
    output [0:0] stall_out,
    input [15:0] tile_id
);
wire [15:0] CB_addr_in_0_O;
wire [31:0] CB_addr_in_0_read_config_data;
wire [7:0] CB_addr_in_0_config_config_addr_in;
wire [15:0] CB_addr_in_1_O;
wire [31:0] CB_addr_in_1_read_config_data;
wire [7:0] CB_addr_in_1_config_config_addr_in;
wire [15:0] CB_chain_data_in_0_O;
wire [31:0] CB_chain_data_in_0_read_config_data;
wire [7:0] CB_chain_data_in_0_config_config_addr_in;
wire [15:0] CB_chain_data_in_1_O;
wire [31:0] CB_chain_data_in_1_read_config_data;
wire [7:0] CB_chain_data_in_1_config_config_addr_in;
wire [15:0] CB_data_in_0_O;
wire [31:0] CB_data_in_0_read_config_data;
wire [7:0] CB_data_in_0_config_config_addr_in;
wire [15:0] CB_data_in_1_O;
wire [31:0] CB_data_in_1_read_config_data;
wire [7:0] CB_data_in_1_config_config_addr_in;
wire [0:0] CB_flush_O;
wire [31:0] CB_flush_read_config_data;
wire [7:0] CB_flush_config_config_addr_in;
wire [0:0] CB_ren_in_0_O;
wire [31:0] CB_ren_in_0_read_config_data;
wire [7:0] CB_ren_in_0_config_config_addr_in;
wire [0:0] CB_ren_in_1_O;
wire [31:0] CB_ren_in_1_read_config_data;
wire [7:0] CB_ren_in_1_config_config_addr_in;
wire [0:0] CB_wen_in_0_O;
wire [31:0] CB_wen_in_0_read_config_data;
wire [7:0] CB_wen_in_0_config_config_addr_in;
wire [0:0] CB_wen_in_1_O;
wire [31:0] CB_wen_in_1_read_config_data;
wire [7:0] CB_wen_in_1_config_config_addr_in;
wire DECODE_FEATURE_0_O;
wire DECODE_FEATURE_1_O;
wire DECODE_FEATURE_10_O;
wire DECODE_FEATURE_11_O;
wire DECODE_FEATURE_12_O;
wire DECODE_FEATURE_13_O;
wire DECODE_FEATURE_14_O;
wire DECODE_FEATURE_15_O;
wire DECODE_FEATURE_2_O;
wire DECODE_FEATURE_3_O;
wire DECODE_FEATURE_4_O;
wire DECODE_FEATURE_5_O;
wire DECODE_FEATURE_6_O;
wire DECODE_FEATURE_7_O;
wire DECODE_FEATURE_8_O;
wire DECODE_FEATURE_9_O;
wire FEATURE_AND_0_out;
wire FEATURE_AND_1_out;
wire FEATURE_AND_10_out;
wire FEATURE_AND_11_out;
wire FEATURE_AND_12_out;
wire FEATURE_AND_13_out;
wire FEATURE_AND_14_out;
wire FEATURE_AND_15_out;
wire FEATURE_AND_2_out;
wire FEATURE_AND_3_out;
wire FEATURE_AND_4_out;
wire FEATURE_AND_5_out;
wire FEATURE_AND_6_out;
wire FEATURE_AND_7_out;
wire FEATURE_AND_8_out;
wire FEATURE_AND_9_out;
wire [15:0] MemCore_inst0_data_out_0;
wire [15:0] MemCore_inst0_data_out_1;
wire [0:0] MemCore_inst0_empty;
wire [0:0] MemCore_inst0_full;
wire [31:0] MemCore_inst0_read_config_data;
wire [31:0] MemCore_inst0_read_config_data_1;
wire [31:0] MemCore_inst0_read_config_data_2;
wire [0:0] MemCore_inst0_sram_ready_out;
wire [0:0] MemCore_inst0_stencil_valid;
wire [0:0] MemCore_inst0_valid_out_0;
wire [0:0] MemCore_inst0_valid_out_1;
wire [7:0] MemCore_inst0_config_1_config_addr_in;
wire [7:0] MemCore_inst0_config_2_config_addr_in;
wire [7:0] MemCore_inst0_config_config_addr_in;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T0_EAST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T0_NORTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T0_SOUTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T0_WEST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T1_EAST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T1_NORTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T1_SOUTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T1_WEST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T2_EAST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T2_NORTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T2_SOUTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T2_WEST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T3_EAST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T3_NORTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T3_SOUTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T3_WEST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T4_EAST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T4_NORTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T4_SOUTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_MemCore_SB_T4_WEST_SB_OUT_B16;
wire [31:0] SB_ID0_5TRACKS_B16_MemCore_read_config_data;
wire [7:0] SB_ID0_5TRACKS_B16_MemCore_config_config_addr_in;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_OUT_B1;
wire [31:0] SB_ID0_5TRACKS_B1_MemCore_read_config_data;
wire [7:0] SB_ID0_5TRACKS_B1_MemCore_config_config_addr_in;
wire [0:0] WIRE_SB_T0_EAST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T0_EAST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T0_NORTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T0_NORTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T0_SOUTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T0_SOUTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T0_WEST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T0_WEST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T1_EAST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T1_EAST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T1_NORTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T1_NORTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T1_SOUTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T1_SOUTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T1_WEST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T1_WEST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T2_EAST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T2_EAST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T2_NORTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T2_NORTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T2_SOUTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T2_SOUTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T2_WEST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T2_WEST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T3_EAST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T3_EAST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T3_NORTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T3_NORTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T3_SOUTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T3_SOUTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T3_WEST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T3_WEST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T4_EAST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T4_EAST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T4_NORTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T4_NORTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T4_SOUTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T4_SOUTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T4_WEST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T4_WEST_SB_IN_B16_O;
wire and_inst0_out;
wire and_inst1_out;
wire [7:0] const_0_8_out;
wire [8:0] const_511_9_out;
wire coreir_eq_16_inst0_out;
wire [31:0] read_config_data_or_inst0_out;
wire [31:0] read_data_mux_O;
wire [7:0] read_data_mux_S_in;
wire [31:0] self_config_config_addr_out;
CB_addr_in_0 CB_addr_in_0 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .O(CB_addr_in_0_O),
    .clk(clk),
    .config_config_addr(CB_addr_in_0_config_config_addr_in),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_3_out),
    .read_config_data(CB_addr_in_0_read_config_data),
    .reset(reset)
);
mantle_wire__typeBitIn8 CB_addr_in_0_config_config_addr (
    .in(CB_addr_in_0_config_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
CB_addr_in_1 CB_addr_in_1 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .O(CB_addr_in_1_O),
    .clk(clk),
    .config_config_addr(CB_addr_in_1_config_config_addr_in),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_4_out),
    .read_config_data(CB_addr_in_1_read_config_data),
    .reset(reset)
);
mantle_wire__typeBitIn8 CB_addr_in_1_config_config_addr (
    .in(CB_addr_in_1_config_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
CB_chain_data_in_0 CB_chain_data_in_0 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .O(CB_chain_data_in_0_O),
    .clk(clk),
    .config_config_addr(CB_chain_data_in_0_config_config_addr_in),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_5_out),
    .read_config_data(CB_chain_data_in_0_read_config_data),
    .reset(reset)
);
mantle_wire__typeBitIn8 CB_chain_data_in_0_config_config_addr (
    .in(CB_chain_data_in_0_config_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
CB_chain_data_in_1 CB_chain_data_in_1 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .O(CB_chain_data_in_1_O),
    .clk(clk),
    .config_config_addr(CB_chain_data_in_1_config_config_addr_in),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_6_out),
    .read_config_data(CB_chain_data_in_1_read_config_data),
    .reset(reset)
);
mantle_wire__typeBitIn8 CB_chain_data_in_1_config_config_addr (
    .in(CB_chain_data_in_1_config_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
CB_data_in_0 CB_data_in_0 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .O(CB_data_in_0_O),
    .clk(clk),
    .config_config_addr(CB_data_in_0_config_config_addr_in),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_7_out),
    .read_config_data(CB_data_in_0_read_config_data),
    .reset(reset)
);
mantle_wire__typeBitIn8 CB_data_in_0_config_config_addr (
    .in(CB_data_in_0_config_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
CB_data_in_1 CB_data_in_1 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .O(CB_data_in_1_O),
    .clk(clk),
    .config_config_addr(CB_data_in_1_config_config_addr_in),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_8_out),
    .read_config_data(CB_data_in_1_read_config_data),
    .reset(reset)
);
mantle_wire__typeBitIn8 CB_data_in_1_config_config_addr (
    .in(CB_data_in_1_config_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
CB_flush CB_flush (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .O(CB_flush_O),
    .clk(clk),
    .config_config_addr(CB_flush_config_config_addr_in),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_9_out),
    .read_config_data(CB_flush_read_config_data),
    .reset(reset)
);
mantle_wire__typeBitIn8 CB_flush_config_config_addr (
    .in(CB_flush_config_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
CB_ren_in_0 CB_ren_in_0 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .O(CB_ren_in_0_O),
    .clk(clk),
    .config_config_addr(CB_ren_in_0_config_config_addr_in),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_10_out),
    .read_config_data(CB_ren_in_0_read_config_data),
    .reset(reset)
);
mantle_wire__typeBitIn8 CB_ren_in_0_config_config_addr (
    .in(CB_ren_in_0_config_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
CB_ren_in_1 CB_ren_in_1 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .O(CB_ren_in_1_O),
    .clk(clk),
    .config_config_addr(CB_ren_in_1_config_config_addr_in),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_11_out),
    .read_config_data(CB_ren_in_1_read_config_data),
    .reset(reset)
);
mantle_wire__typeBitIn8 CB_ren_in_1_config_config_addr (
    .in(CB_ren_in_1_config_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
CB_wen_in_0 CB_wen_in_0 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .O(CB_wen_in_0_O),
    .clk(clk),
    .config_config_addr(CB_wen_in_0_config_config_addr_in),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_12_out),
    .read_config_data(CB_wen_in_0_read_config_data),
    .reset(reset)
);
mantle_wire__typeBitIn8 CB_wen_in_0_config_config_addr (
    .in(CB_wen_in_0_config_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
CB_wen_in_1 CB_wen_in_1 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .O(CB_wen_in_1_O),
    .clk(clk),
    .config_config_addr(CB_wen_in_1_config_config_addr_in),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_13_out),
    .read_config_data(CB_wen_in_1_read_config_data),
    .reset(reset)
);
mantle_wire__typeBitIn8 CB_wen_in_1_config_config_addr (
    .in(CB_wen_in_1_config_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
Decode08 DECODE_FEATURE_0 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_0_O)
);
Decode18 DECODE_FEATURE_1 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_1_O)
);
Decode108 DECODE_FEATURE_10 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_10_O)
);
Decode118 DECODE_FEATURE_11 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_11_O)
);
Decode128 DECODE_FEATURE_12 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_12_O)
);
Decode138 DECODE_FEATURE_13 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_13_O)
);
Decode148 DECODE_FEATURE_14 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_14_O)
);
Decode158 DECODE_FEATURE_15 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_15_O)
);
Decode28 DECODE_FEATURE_2 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_2_O)
);
Decode38 DECODE_FEATURE_3 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_3_O)
);
Decode48 DECODE_FEATURE_4 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_4_O)
);
Decode58 DECODE_FEATURE_5 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_5_O)
);
Decode68 DECODE_FEATURE_6 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_6_O)
);
Decode78 DECODE_FEATURE_7 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_7_O)
);
Decode88 DECODE_FEATURE_8 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_8_O)
);
Decode98 DECODE_FEATURE_9 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_9_O)
);
corebit_and FEATURE_AND_0 (
    .in0(DECODE_FEATURE_0_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_0_out)
);
corebit_and FEATURE_AND_1 (
    .in0(DECODE_FEATURE_1_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_1_out)
);
corebit_and FEATURE_AND_10 (
    .in0(DECODE_FEATURE_10_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_10_out)
);
corebit_and FEATURE_AND_11 (
    .in0(DECODE_FEATURE_11_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_11_out)
);
corebit_and FEATURE_AND_12 (
    .in0(DECODE_FEATURE_12_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_12_out)
);
corebit_and FEATURE_AND_13 (
    .in0(DECODE_FEATURE_13_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_13_out)
);
corebit_and FEATURE_AND_14 (
    .in0(DECODE_FEATURE_14_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_14_out)
);
corebit_and FEATURE_AND_15 (
    .in0(DECODE_FEATURE_15_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_15_out)
);
corebit_and FEATURE_AND_2 (
    .in0(DECODE_FEATURE_2_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_2_out)
);
corebit_and FEATURE_AND_3 (
    .in0(DECODE_FEATURE_3_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_3_out)
);
corebit_and FEATURE_AND_4 (
    .in0(DECODE_FEATURE_4_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_4_out)
);
corebit_and FEATURE_AND_5 (
    .in0(DECODE_FEATURE_5_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_5_out)
);
corebit_and FEATURE_AND_6 (
    .in0(DECODE_FEATURE_6_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_6_out)
);
corebit_and FEATURE_AND_7 (
    .in0(DECODE_FEATURE_7_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_7_out)
);
corebit_and FEATURE_AND_8 (
    .in0(DECODE_FEATURE_8_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_8_out)
);
corebit_and FEATURE_AND_9 (
    .in0(DECODE_FEATURE_9_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_9_out)
);
MemCore MemCore_inst0 (
    .addr_in_0(CB_addr_in_0_O),
    .addr_in_1(CB_addr_in_1_O),
    .chain_data_in_0(CB_chain_data_in_0_O),
    .chain_data_in_1(CB_chain_data_in_1_O),
    .clk(clk),
    .config_1_config_addr(MemCore_inst0_config_1_config_addr_in),
    .config_1_config_data(config_config_data),
    .config_1_read(config_read),
    .config_1_write(FEATURE_AND_1_out),
    .config_2_config_addr(MemCore_inst0_config_2_config_addr_in),
    .config_2_config_data(config_config_data),
    .config_2_read(config_read),
    .config_2_write(FEATURE_AND_2_out),
    .config_config_addr(MemCore_inst0_config_config_addr_in),
    .config_config_data(config_config_data),
    .config_en_0(DECODE_FEATURE_1_O),
    .config_en_1(DECODE_FEATURE_2_O),
    .config_read(config_read),
    .config_write(FEATURE_AND_0_out),
    .data_in_0(CB_data_in_0_O),
    .data_in_1(CB_data_in_1_O),
    .data_out_0(MemCore_inst0_data_out_0),
    .data_out_1(MemCore_inst0_data_out_1),
    .empty(MemCore_inst0_empty),
    .flush(CB_flush_O),
    .full(MemCore_inst0_full),
    .read_config_data(MemCore_inst0_read_config_data),
    .read_config_data_1(MemCore_inst0_read_config_data_1),
    .read_config_data_2(MemCore_inst0_read_config_data_2),
    .ren_in_0(CB_ren_in_0_O),
    .ren_in_1(CB_ren_in_1_O),
    .reset(reset),
    .sram_ready_out(MemCore_inst0_sram_ready_out),
    .stall(stall),
    .stencil_valid(MemCore_inst0_stencil_valid),
    .valid_out_0(MemCore_inst0_valid_out_0),
    .valid_out_1(MemCore_inst0_valid_out_1),
    .wen_in_0(CB_wen_in_0_O),
    .wen_in_1(CB_wen_in_1_O)
);
mantle_wire__typeBitIn8 MemCore_inst0_config_1_config_addr (
    .in(MemCore_inst0_config_1_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
mantle_wire__typeBitIn8 MemCore_inst0_config_2_config_addr (
    .in(MemCore_inst0_config_2_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
mantle_wire__typeBitIn8 MemCore_inst0_config_config_addr (
    .in(MemCore_inst0_config_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
SB_ID0_5TRACKS_B16_MemCore SB_ID0_5TRACKS_B16_MemCore (
    .SB_T0_EAST_SB_IN_B16(SB_T0_EAST_SB_IN_B16),
    .SB_T0_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B16(SB_T0_NORTH_SB_IN_B16),
    .SB_T0_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B16(SB_T0_SOUTH_SB_IN_B16),
    .SB_T0_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B16(SB_T0_WEST_SB_IN_B16),
    .SB_T0_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B16(SB_T1_EAST_SB_IN_B16),
    .SB_T1_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B16(SB_T1_NORTH_SB_IN_B16),
    .SB_T1_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B16(SB_T1_SOUTH_SB_IN_B16),
    .SB_T1_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B16(SB_T1_WEST_SB_IN_B16),
    .SB_T1_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B16(SB_T2_EAST_SB_IN_B16),
    .SB_T2_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B16(SB_T2_NORTH_SB_IN_B16),
    .SB_T2_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B16(SB_T2_SOUTH_SB_IN_B16),
    .SB_T2_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B16(SB_T2_WEST_SB_IN_B16),
    .SB_T2_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B16(SB_T3_EAST_SB_IN_B16),
    .SB_T3_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B16(SB_T3_NORTH_SB_IN_B16),
    .SB_T3_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B16(SB_T3_SOUTH_SB_IN_B16),
    .SB_T3_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B16(SB_T3_WEST_SB_IN_B16),
    .SB_T3_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B16(SB_T4_EAST_SB_IN_B16),
    .SB_T4_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B16(SB_T4_NORTH_SB_IN_B16),
    .SB_T4_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B16(SB_T4_SOUTH_SB_IN_B16),
    .SB_T4_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B16(SB_T4_WEST_SB_IN_B16),
    .SB_T4_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_MemCore_SB_T4_WEST_SB_OUT_B16),
    .clk(clk),
    .config_config_addr(SB_ID0_5TRACKS_B16_MemCore_config_config_addr_in),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_15_out),
    .data_out_0(MemCore_inst0_data_out_0),
    .data_out_1(MemCore_inst0_data_out_1),
    .read_config_data(SB_ID0_5TRACKS_B16_MemCore_read_config_data),
    .reset(reset),
    .stall(stall)
);
mantle_wire__typeBitIn8 SB_ID0_5TRACKS_B16_MemCore_config_config_addr (
    .in(SB_ID0_5TRACKS_B16_MemCore_config_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
SB_ID0_5TRACKS_B1_MemCore SB_ID0_5TRACKS_B1_MemCore (
    .SB_T0_EAST_SB_IN_B1(SB_T0_EAST_SB_IN_B1),
    .SB_T0_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B1(SB_T0_NORTH_SB_IN_B1),
    .SB_T0_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B1(SB_T0_SOUTH_SB_IN_B1),
    .SB_T0_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B1(SB_T0_WEST_SB_IN_B1),
    .SB_T0_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B1(SB_T1_EAST_SB_IN_B1),
    .SB_T1_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B1(SB_T1_NORTH_SB_IN_B1),
    .SB_T1_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B1(SB_T1_SOUTH_SB_IN_B1),
    .SB_T1_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B1(SB_T1_WEST_SB_IN_B1),
    .SB_T1_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B1(SB_T2_EAST_SB_IN_B1),
    .SB_T2_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B1(SB_T2_NORTH_SB_IN_B1),
    .SB_T2_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B1(SB_T2_SOUTH_SB_IN_B1),
    .SB_T2_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B1(SB_T2_WEST_SB_IN_B1),
    .SB_T2_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B1(SB_T3_EAST_SB_IN_B1),
    .SB_T3_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B1(SB_T3_NORTH_SB_IN_B1),
    .SB_T3_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B1(SB_T3_SOUTH_SB_IN_B1),
    .SB_T3_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B1(SB_T3_WEST_SB_IN_B1),
    .SB_T3_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B1(SB_T4_EAST_SB_IN_B1),
    .SB_T4_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B1(SB_T4_NORTH_SB_IN_B1),
    .SB_T4_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B1(SB_T4_SOUTH_SB_IN_B1),
    .SB_T4_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B1(SB_T4_WEST_SB_IN_B1),
    .SB_T4_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_OUT_B1),
    .clk(clk),
    .config_config_addr(SB_ID0_5TRACKS_B1_MemCore_config_config_addr_in),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_14_out),
    .empty(MemCore_inst0_empty),
    .full(MemCore_inst0_full),
    .read_config_data(SB_ID0_5TRACKS_B1_MemCore_read_config_data),
    .reset(reset),
    .sram_ready_out(MemCore_inst0_sram_ready_out),
    .stall(stall),
    .stencil_valid(MemCore_inst0_stencil_valid),
    .valid_out_0(MemCore_inst0_valid_out_0),
    .valid_out_1(MemCore_inst0_valid_out_1)
);
mantle_wire__typeBitIn8 SB_ID0_5TRACKS_B1_MemCore_config_config_addr (
    .in(SB_ID0_5TRACKS_B1_MemCore_config_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
MuxWrapper_1_1 WIRE_SB_T0_EAST_SB_IN_B1 (
    .I(SB_T0_EAST_SB_IN_B1),
    .O(WIRE_SB_T0_EAST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T0_EAST_SB_IN_B16 (
    .I(SB_T0_EAST_SB_IN_B16),
    .O(WIRE_SB_T0_EAST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T0_NORTH_SB_IN_B1 (
    .I(SB_T0_NORTH_SB_IN_B1),
    .O(WIRE_SB_T0_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T0_NORTH_SB_IN_B16 (
    .I(SB_T0_NORTH_SB_IN_B16),
    .O(WIRE_SB_T0_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T0_SOUTH_SB_IN_B1 (
    .I(SB_T0_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T0_SOUTH_SB_IN_B16 (
    .I(SB_T0_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T0_WEST_SB_IN_B1 (
    .I(SB_T0_WEST_SB_IN_B1),
    .O(WIRE_SB_T0_WEST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T0_WEST_SB_IN_B16 (
    .I(SB_T0_WEST_SB_IN_B16),
    .O(WIRE_SB_T0_WEST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T1_EAST_SB_IN_B1 (
    .I(SB_T1_EAST_SB_IN_B1),
    .O(WIRE_SB_T1_EAST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T1_EAST_SB_IN_B16 (
    .I(SB_T1_EAST_SB_IN_B16),
    .O(WIRE_SB_T1_EAST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T1_NORTH_SB_IN_B1 (
    .I(SB_T1_NORTH_SB_IN_B1),
    .O(WIRE_SB_T1_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T1_NORTH_SB_IN_B16 (
    .I(SB_T1_NORTH_SB_IN_B16),
    .O(WIRE_SB_T1_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T1_SOUTH_SB_IN_B1 (
    .I(SB_T1_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T1_SOUTH_SB_IN_B16 (
    .I(SB_T1_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T1_WEST_SB_IN_B1 (
    .I(SB_T1_WEST_SB_IN_B1),
    .O(WIRE_SB_T1_WEST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T1_WEST_SB_IN_B16 (
    .I(SB_T1_WEST_SB_IN_B16),
    .O(WIRE_SB_T1_WEST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T2_EAST_SB_IN_B1 (
    .I(SB_T2_EAST_SB_IN_B1),
    .O(WIRE_SB_T2_EAST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T2_EAST_SB_IN_B16 (
    .I(SB_T2_EAST_SB_IN_B16),
    .O(WIRE_SB_T2_EAST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T2_NORTH_SB_IN_B1 (
    .I(SB_T2_NORTH_SB_IN_B1),
    .O(WIRE_SB_T2_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T2_NORTH_SB_IN_B16 (
    .I(SB_T2_NORTH_SB_IN_B16),
    .O(WIRE_SB_T2_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T2_SOUTH_SB_IN_B1 (
    .I(SB_T2_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T2_SOUTH_SB_IN_B16 (
    .I(SB_T2_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T2_WEST_SB_IN_B1 (
    .I(SB_T2_WEST_SB_IN_B1),
    .O(WIRE_SB_T2_WEST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T2_WEST_SB_IN_B16 (
    .I(SB_T2_WEST_SB_IN_B16),
    .O(WIRE_SB_T2_WEST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T3_EAST_SB_IN_B1 (
    .I(SB_T3_EAST_SB_IN_B1),
    .O(WIRE_SB_T3_EAST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T3_EAST_SB_IN_B16 (
    .I(SB_T3_EAST_SB_IN_B16),
    .O(WIRE_SB_T3_EAST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T3_NORTH_SB_IN_B1 (
    .I(SB_T3_NORTH_SB_IN_B1),
    .O(WIRE_SB_T3_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T3_NORTH_SB_IN_B16 (
    .I(SB_T3_NORTH_SB_IN_B16),
    .O(WIRE_SB_T3_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T3_SOUTH_SB_IN_B1 (
    .I(SB_T3_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T3_SOUTH_SB_IN_B16 (
    .I(SB_T3_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T3_WEST_SB_IN_B1 (
    .I(SB_T3_WEST_SB_IN_B1),
    .O(WIRE_SB_T3_WEST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T3_WEST_SB_IN_B16 (
    .I(SB_T3_WEST_SB_IN_B16),
    .O(WIRE_SB_T3_WEST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T4_EAST_SB_IN_B1 (
    .I(SB_T4_EAST_SB_IN_B1),
    .O(WIRE_SB_T4_EAST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T4_EAST_SB_IN_B16 (
    .I(SB_T4_EAST_SB_IN_B16),
    .O(WIRE_SB_T4_EAST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T4_NORTH_SB_IN_B1 (
    .I(SB_T4_NORTH_SB_IN_B1),
    .O(WIRE_SB_T4_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T4_NORTH_SB_IN_B16 (
    .I(SB_T4_NORTH_SB_IN_B16),
    .O(WIRE_SB_T4_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T4_SOUTH_SB_IN_B1 (
    .I(SB_T4_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T4_SOUTH_SB_IN_B16 (
    .I(SB_T4_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T4_WEST_SB_IN_B1 (
    .I(SB_T4_WEST_SB_IN_B1),
    .O(WIRE_SB_T4_WEST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T4_WEST_SB_IN_B16 (
    .I(SB_T4_WEST_SB_IN_B16),
    .O(WIRE_SB_T4_WEST_SB_IN_B16_O)
);
corebit_and and_inst0 (
    .in0(coreir_eq_16_inst0_out),
    .in1(config_read[0]),
    .out(and_inst0_out)
);
corebit_and and_inst1 (
    .in0(coreir_eq_16_inst0_out),
    .in1(config_write[0]),
    .out(and_inst1_out)
);
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
coreir_const #(
    .value(9'h1ff),
    .width(9)
) const_511_9 (
    .out(const_511_9_out)
);
coreir_eq #(
    .width(16)
) coreir_eq_16_inst0 (
    .in0(tile_id),
    .in1(self_config_config_addr_out[15:0]),
    .out(coreir_eq_16_inst0_out)
);
coreir_or #(
    .width(32)
) read_config_data_or_inst0 (
    .in0(read_data_mux_O),
    .in1(read_config_data_in),
    .out(read_config_data_or_inst0_out)
);
MuxWithDefaultWrapper_16_32_8_0 read_data_mux (
    .EN(and_inst0_out),
    .I_0(MemCore_inst0_read_config_data),
    .I_1(MemCore_inst0_read_config_data_1),
    .I_10(CB_ren_in_0_read_config_data),
    .I_11(CB_ren_in_1_read_config_data),
    .I_12(CB_wen_in_0_read_config_data),
    .I_13(CB_wen_in_1_read_config_data),
    .I_14(SB_ID0_5TRACKS_B1_MemCore_read_config_data),
    .I_15(SB_ID0_5TRACKS_B16_MemCore_read_config_data),
    .I_2(MemCore_inst0_read_config_data_2),
    .I_3(CB_addr_in_0_read_config_data),
    .I_4(CB_addr_in_1_read_config_data),
    .I_5(CB_chain_data_in_0_read_config_data),
    .I_6(CB_chain_data_in_1_read_config_data),
    .I_7(CB_data_in_0_read_config_data),
    .I_8(CB_data_in_1_read_config_data),
    .I_9(CB_flush_read_config_data),
    .O(read_data_mux_O),
    .S(read_data_mux_S_in)
);
mantle_wire__typeBitIn8 read_data_mux_S (
    .in(read_data_mux_S_in),
    .out(self_config_config_addr_out[23:16])
);
mantle_wire__typeBit32 self_config_config_addr (
    .in(config_config_addr),
    .out(self_config_config_addr_out)
);
assign SB_T0_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T0_EAST_SB_OUT_B1;
assign SB_T0_EAST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T0_EAST_SB_OUT_B16;
assign SB_T0_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T0_NORTH_SB_OUT_B1;
assign SB_T0_NORTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T0_NORTH_SB_OUT_B16;
assign SB_T0_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T0_SOUTH_SB_OUT_B1;
assign SB_T0_SOUTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T0_SOUTH_SB_OUT_B16;
assign SB_T0_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T0_WEST_SB_OUT_B1;
assign SB_T0_WEST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T0_WEST_SB_OUT_B16;
assign SB_T1_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T1_EAST_SB_OUT_B1;
assign SB_T1_EAST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T1_EAST_SB_OUT_B16;
assign SB_T1_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T1_NORTH_SB_OUT_B1;
assign SB_T1_NORTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T1_NORTH_SB_OUT_B16;
assign SB_T1_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T1_SOUTH_SB_OUT_B1;
assign SB_T1_SOUTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T1_SOUTH_SB_OUT_B16;
assign SB_T1_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T1_WEST_SB_OUT_B1;
assign SB_T1_WEST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T1_WEST_SB_OUT_B16;
assign SB_T2_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T2_EAST_SB_OUT_B1;
assign SB_T2_EAST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T2_EAST_SB_OUT_B16;
assign SB_T2_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T2_NORTH_SB_OUT_B1;
assign SB_T2_NORTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T2_NORTH_SB_OUT_B16;
assign SB_T2_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T2_SOUTH_SB_OUT_B1;
assign SB_T2_SOUTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T2_SOUTH_SB_OUT_B16;
assign SB_T2_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T2_WEST_SB_OUT_B1;
assign SB_T2_WEST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T2_WEST_SB_OUT_B16;
assign SB_T3_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T3_EAST_SB_OUT_B1;
assign SB_T3_EAST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T3_EAST_SB_OUT_B16;
assign SB_T3_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T3_NORTH_SB_OUT_B1;
assign SB_T3_NORTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T3_NORTH_SB_OUT_B16;
assign SB_T3_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T3_SOUTH_SB_OUT_B1;
assign SB_T3_SOUTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T3_SOUTH_SB_OUT_B16;
assign SB_T3_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T3_WEST_SB_OUT_B1;
assign SB_T3_WEST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T3_WEST_SB_OUT_B16;
assign SB_T4_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T4_EAST_SB_OUT_B1;
assign SB_T4_EAST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T4_EAST_SB_OUT_B16;
assign SB_T4_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T4_NORTH_SB_OUT_B1;
assign SB_T4_NORTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T4_NORTH_SB_OUT_B16;
assign SB_T4_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T4_SOUTH_SB_OUT_B1;
assign SB_T4_SOUTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T4_SOUTH_SB_OUT_B16;
assign SB_T4_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_MemCore_SB_T4_WEST_SB_OUT_B1;
assign SB_T4_WEST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_MemCore_SB_T4_WEST_SB_OUT_B16;
assign clk_out = clk;
assign config_out_config_addr = config_config_addr;
assign config_out_config_data = config_config_data;
assign config_out_read = config_read;
assign config_out_write = config_write;
assign hi = const_511_9_out;
assign lo = const_0_8_out;
assign read_config_data = read_config_data_or_inst0_out;
assign reset_out = reset;
assign stall_out = stall;
endmodule

module BIT_ALU (
    input [1:0] alu,
    input [15:0] a,
    input [15:0] b,
    output [15:0] O0,
    output O1,
    output O2,
    output O3,
    output O4,
    output O5,
    input CLK,
    input ASYNCRESET
);
wire [0:0] Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out;
wire [15:0] Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out;
wire bit_const_0_None_out;
wire [15:0] const_0_16_out;
wire [1:0] const_0_2_out;
wire [1:0] const_1_2_out;
wire [15:0] magma_Bits_16_and_inst0_out;
wire magma_Bits_16_eq_inst0_out;
wire [15:0] magma_Bits_16_or_inst0_out;
wire [15:0] magma_Bits_16_xor_inst0_out;
wire magma_Bits_2_eq_inst0_out;
wire magma_Bits_2_eq_inst1_out;
coreir_mux #(
    .width(1)
) Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(bit_const_0_None_out),
    .in1(bit_const_0_None_out),
    .sel(magma_Bits_2_eq_inst0_out),
    .out(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(bit_const_0_None_out),
    .sel(magma_Bits_2_eq_inst1_out),
    .out(Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(magma_Bits_16_xor_inst0_out),
    .in1(magma_Bits_16_or_inst0_out),
    .sel(magma_Bits_2_eq_inst0_out),
    .out(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(magma_Bits_16_and_inst0_out),
    .sel(magma_Bits_2_eq_inst1_out),
    .out(Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out)
);
corebit_const #(
    .value(1'b0)
) bit_const_0_None (
    .out(bit_const_0_None_out)
);
coreir_const #(
    .value(16'h0000),
    .width(16)
) const_0_16 (
    .out(const_0_16_out)
);
coreir_const #(
    .value(2'h0),
    .width(2)
) const_0_2 (
    .out(const_0_2_out)
);
coreir_const #(
    .value(2'h1),
    .width(2)
) const_1_2 (
    .out(const_1_2_out)
);
coreir_and #(
    .width(16)
) magma_Bits_16_and_inst0 (
    .in0(a),
    .in1(b),
    .out(magma_Bits_16_and_inst0_out)
);
coreir_eq #(
    .width(16)
) magma_Bits_16_eq_inst0 (
    .in0(Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(const_0_16_out),
    .out(magma_Bits_16_eq_inst0_out)
);
coreir_or #(
    .width(16)
) magma_Bits_16_or_inst0 (
    .in0(a),
    .in1(b),
    .out(magma_Bits_16_or_inst0_out)
);
coreir_xor #(
    .width(16)
) magma_Bits_16_xor_inst0 (
    .in0(a),
    .in1(b),
    .out(magma_Bits_16_xor_inst0_out)
);
coreir_eq #(
    .width(2)
) magma_Bits_2_eq_inst0 (
    .in0(alu),
    .in1(const_0_2_out),
    .out(magma_Bits_2_eq_inst0_out)
);
coreir_eq #(
    .width(2)
) magma_Bits_2_eq_inst1 (
    .in0(alu),
    .in1(const_1_2_out),
    .out(magma_Bits_2_eq_inst1_out)
);
assign O0 = Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out;
assign O1 = Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out[0];
assign O2 = magma_Bits_16_eq_inst0_out;
assign O3 = Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out[15];
assign O4 = bit_const_0_None_out;
assign O5 = bit_const_0_None_out;
endmodule

module ADD (
    input [15:0] a,
    input [15:0] b,
    output [15:0] O0,
    output O1,
    output O2,
    output O3,
    output O4,
    output O5,
    input CLK,
    input ASYNCRESET
);
wire bit_const_0_None_out;
wire [15:0] const_0_16_out;
wire [16:0] const_0_17_out;
wire magma_Bit_and_inst0_out;
wire magma_Bit_and_inst1_out;
wire magma_Bit_and_inst2_out;
wire magma_Bit_and_inst3_out;
wire magma_Bit_not_inst0_out;
wire magma_Bit_not_inst1_out;
wire magma_Bit_not_inst2_out;
wire magma_Bit_or_inst0_out;
wire magma_Bits_16_eq_inst0_out;
wire [16:0] magma_Bits_17_add_inst0_out;
wire [16:0] magma_Bits_17_add_inst1_out;
corebit_const #(
    .value(1'b0)
) bit_const_0_None (
    .out(bit_const_0_None_out)
);
coreir_const #(
    .value(16'h0000),
    .width(16)
) const_0_16 (
    .out(const_0_16_out)
);
coreir_const #(
    .value(17'h00000),
    .width(17)
) const_0_17 (
    .out(const_0_17_out)
);
corebit_and magma_Bit_and_inst0 (
    .in0(a[15]),
    .in1(b[15]),
    .out(magma_Bit_and_inst0_out)
);
corebit_and magma_Bit_and_inst1 (
    .in0(magma_Bit_and_inst0_out),
    .in1(magma_Bit_not_inst0_out),
    .out(magma_Bit_and_inst1_out)
);
corebit_and magma_Bit_and_inst2 (
    .in0(magma_Bit_not_inst1_out),
    .in1(magma_Bit_not_inst2_out),
    .out(magma_Bit_and_inst2_out)
);
corebit_and magma_Bit_and_inst3 (
    .in0(magma_Bit_and_inst2_out),
    .in1(magma_Bits_17_add_inst1_out[15]),
    .out(magma_Bit_and_inst3_out)
);
corebit_not magma_Bit_not_inst0 (
    .in(magma_Bits_17_add_inst1_out[15]),
    .out(magma_Bit_not_inst0_out)
);
corebit_not magma_Bit_not_inst1 (
    .in(a[15]),
    .out(magma_Bit_not_inst1_out)
);
corebit_not magma_Bit_not_inst2 (
    .in(b[15]),
    .out(magma_Bit_not_inst2_out)
);
corebit_or magma_Bit_or_inst0 (
    .in0(magma_Bit_and_inst1_out),
    .in1(magma_Bit_and_inst3_out),
    .out(magma_Bit_or_inst0_out)
);
coreir_eq #(
    .width(16)
) magma_Bits_16_eq_inst0 (
    .in0(magma_Bits_17_add_inst1_out[15:0]),
    .in1(const_0_16_out),
    .out(magma_Bits_16_eq_inst0_out)
);
wire [16:0] magma_Bits_17_add_inst0_in0;
assign magma_Bits_17_add_inst0_in0 = {bit_const_0_None_out,a[15:0]};
wire [16:0] magma_Bits_17_add_inst0_in1;
assign magma_Bits_17_add_inst0_in1 = {bit_const_0_None_out,b[15:0]};
coreir_add #(
    .width(17)
) magma_Bits_17_add_inst0 (
    .in0(magma_Bits_17_add_inst0_in0),
    .in1(magma_Bits_17_add_inst0_in1),
    .out(magma_Bits_17_add_inst0_out)
);
coreir_add #(
    .width(17)
) magma_Bits_17_add_inst1 (
    .in0(magma_Bits_17_add_inst0_out),
    .in1(const_0_17_out),
    .out(magma_Bits_17_add_inst1_out)
);
assign O0 = magma_Bits_17_add_inst1_out[15:0];
assign O1 = magma_Bits_17_add_inst1_out[16];
assign O2 = magma_Bits_16_eq_inst0_out;
assign O3 = magma_Bits_17_add_inst1_out[15];
assign O4 = magma_Bits_17_add_inst1_out[16];
assign O5 = magma_Bit_or_inst0_out;
endmodule

module ABSD (
    input [15:0] a,
    input [15:0] b,
    output [15:0] O0,
    output O1,
    output O2,
    output O3,
    output O4,
    output O5,
    input CLK,
    input ASYNCRESET
);
wire [15:0] Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst0_I0_in;
wire bit_const_0_None_out;
wire [15:0] const_0_16_out;
wire [16:0] const_1_17_out;
wire magma_Bits_16_eq_inst0_out;
wire [15:0] magma_Bits_16_neg_inst0_out;
wire [15:0] magma_Bits_16_not_inst0_out;
wire magma_Bits_16_slt_inst0_out;
wire [16:0] magma_Bits_17_add_inst0_out;
wire [16:0] magma_Bits_17_add_inst1_out;
coreir_mux #(
    .width(16)
) Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst0_I0_in),
    .in1(magma_Bits_16_neg_inst0_out),
    .sel(magma_Bits_16_slt_inst0_out),
    .out(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
mantle_wire__typeBitIn16 Mux2xBits16_inst0_I0 (
    .in(Mux2xBits16_inst0_I0_in),
    .out(magma_Bits_17_add_inst1_out[15:0])
);
corebit_const #(
    .value(1'b0)
) bit_const_0_None (
    .out(bit_const_0_None_out)
);
coreir_const #(
    .value(16'h0000),
    .width(16)
) const_0_16 (
    .out(const_0_16_out)
);
coreir_const #(
    .value(17'h00001),
    .width(17)
) const_1_17 (
    .out(const_1_17_out)
);
coreir_eq #(
    .width(16)
) magma_Bits_16_eq_inst0 (
    .in0(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(const_0_16_out),
    .out(magma_Bits_16_eq_inst0_out)
);
coreir_neg #(
    .width(16)
) magma_Bits_16_neg_inst0 (
    .in(magma_Bits_17_add_inst1_out[15:0]),
    .out(magma_Bits_16_neg_inst0_out)
);
coreir_not #(
    .width(16)
) magma_Bits_16_not_inst0 (
    .in(b),
    .out(magma_Bits_16_not_inst0_out)
);
coreir_slt #(
    .width(16)
) magma_Bits_16_slt_inst0 (
    .in0(magma_Bits_17_add_inst1_out[15:0]),
    .in1(const_0_16_out),
    .out(magma_Bits_16_slt_inst0_out)
);
wire [16:0] magma_Bits_17_add_inst0_in0;
assign magma_Bits_17_add_inst0_in0 = {bit_const_0_None_out,a[15:0]};
wire [16:0] magma_Bits_17_add_inst0_in1;
assign magma_Bits_17_add_inst0_in1 = {bit_const_0_None_out,magma_Bits_16_not_inst0_out[15:0]};
coreir_add #(
    .width(17)
) magma_Bits_17_add_inst0 (
    .in0(magma_Bits_17_add_inst0_in0),
    .in1(magma_Bits_17_add_inst0_in1),
    .out(magma_Bits_17_add_inst0_out)
);
coreir_add #(
    .width(17)
) magma_Bits_17_add_inst1 (
    .in0(magma_Bits_17_add_inst0_out),
    .in1(const_1_17_out),
    .out(magma_Bits_17_add_inst1_out)
);
assign O0 = Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
assign O1 = bit_const_0_None_out;
assign O2 = magma_Bits_16_eq_inst0_out;
assign O3 = Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out[15];
assign O4 = bit_const_0_None_out;
assign O5 = bit_const_0_None_out;
endmodule

module PE_gen (
    input [56:0] inst,
    input [50:0] inputs,
    input clk_en,
    output [16:0] O,
    input CLK,
    input ASYNCRESET
);
wire [15:0] ABSD_inst0_O0;
wire ABSD_inst0_O1;
wire ABSD_inst0_O2;
wire ABSD_inst0_O3;
wire ABSD_inst0_O4;
wire ABSD_inst0_O5;
wire [15:0] ADD_inst0_O0;
wire ADD_inst0_O1;
wire ADD_inst0_O2;
wire ADD_inst0_O3;
wire ADD_inst0_O4;
wire ADD_inst0_O5;
wire [15:0] ADD_inst1_O0;
wire ADD_inst1_O1;
wire ADD_inst1_O2;
wire ADD_inst1_O3;
wire ADD_inst1_O4;
wire ADD_inst1_O5;
wire [15:0] BIT_ALU_inst0_O0;
wire BIT_ALU_inst0_O1;
wire BIT_ALU_inst0_O2;
wire BIT_ALU_inst0_O3;
wire BIT_ALU_inst0_O4;
wire BIT_ALU_inst0_O5;
wire Cond_inst0_O;
wire Cond_inst1_O;
wire Cond_inst2_O;
wire [15:0] GTE_inst0_O0;
wire GTE_inst0_O1;
wire GTE_inst0_O2;
wire GTE_inst0_O3;
wire GTE_inst0_O4;
wire GTE_inst0_O5;
wire [15:0] LTE_inst0_O0;
wire LTE_inst0_O1;
wire LTE_inst0_O2;
wire LTE_inst0_O3;
wire LTE_inst0_O4;
wire LTE_inst0_O5;
wire LUT_inst0_O;
wire [15:0] MUL_inst0_O;
wire [0:0] Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out;
wire [0:0] Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out;
wire [15:0] Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst0_I0_in;
wire [15:0] Mux2xBits16_inst0_I1_in;
wire [15:0] Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst10$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst11$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst12$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst13$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst14$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst14_O_out;
wire [15:0] Mux2xBits16_inst1_I1_in;
wire [15:0] Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst2_I0_in;
wire [15:0] Mux2xBits16_inst2_I1_in;
wire [15:0] Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst5$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst6$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst8$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst9$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux2xBits16_inst9_I1_in;
wire [15:0] Mux_inst0$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out;
wire [15:0] Mux_inst0_a_in;
wire [15:0] Mux_inst0_b_in;
wire [15:0] SHR_inst0_O0;
wire SHR_inst0_O1;
wire SHR_inst0_O2;
wire SHR_inst0_O3;
wire SHR_inst0_O4;
wire SHR_inst0_O5;
wire [15:0] SUB_inst0_O0;
wire SUB_inst0_O1;
wire SUB_inst0_O2;
wire SUB_inst0_O3;
wire SUB_inst0_O4;
wire SUB_inst0_O5;
wire [0:0] const_0_1_out;
wire [2:0] const_0_3_out;
wire [3:0] const_0_4_out;
wire [3:0] const_10_4_out;
wire [0:0] const_1_1_out;
wire [2:0] const_1_3_out;
wire [3:0] const_1_4_out;
wire [2:0] const_2_3_out;
wire [3:0] const_2_4_out;
wire [2:0] const_3_3_out;
wire [3:0] const_3_4_out;
wire [2:0] const_4_3_out;
wire [3:0] const_4_4_out;
wire [3:0] const_5_4_out;
wire [3:0] const_6_4_out;
wire [3:0] const_7_4_out;
wire [3:0] const_8_4_out;
wire [3:0] const_9_4_out;
wire magma_Bits_1_eq_inst0_out;
wire magma_Bits_1_eq_inst1_out;
wire magma_Bits_1_eq_inst2_out;
wire magma_Bits_1_eq_inst3_out;
wire magma_Bits_3_eq_inst0_out;
wire magma_Bits_3_eq_inst1_out;
wire magma_Bits_3_eq_inst2_out;
wire magma_Bits_3_eq_inst3_out;
wire magma_Bits_3_eq_inst4_out;
wire magma_Bits_4_eq_inst0_out;
wire magma_Bits_4_eq_inst1_out;
wire magma_Bits_4_eq_inst10_out;
wire magma_Bits_4_eq_inst2_out;
wire magma_Bits_4_eq_inst3_out;
wire magma_Bits_4_eq_inst4_out;
wire magma_Bits_4_eq_inst5_out;
wire magma_Bits_4_eq_inst6_out;
wire magma_Bits_4_eq_inst7_out;
wire magma_Bits_4_eq_inst8_out;
wire magma_Bits_4_eq_inst9_out;
ABSD ABSD_inst0 (
    .a(inputs[47:32]),
    .b(inputs[15:0]),
    .O0(ABSD_inst0_O0),
    .O1(ABSD_inst0_O1),
    .O2(ABSD_inst0_O2),
    .O3(ABSD_inst0_O3),
    .O4(ABSD_inst0_O4),
    .O5(ABSD_inst0_O5),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
ADD ADD_inst0 (
    .a(inputs[15:0]),
    .b(inputs[31:16]),
    .O0(ADD_inst0_O0),
    .O1(ADD_inst0_O1),
    .O2(ADD_inst0_O2),
    .O3(ADD_inst0_O3),
    .O4(ADD_inst0_O4),
    .O5(ADD_inst0_O5),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
ADD ADD_inst1 (
    .a(inputs[47:32]),
    .b(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out),
    .O0(ADD_inst1_O0),
    .O1(ADD_inst1_O1),
    .O2(ADD_inst1_O2),
    .O3(ADD_inst1_O3),
    .O4(ADD_inst1_O4),
    .O5(ADD_inst1_O5),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
BIT_ALU BIT_ALU_inst0 (
    .alu(inst[1:0]),
    .a(inputs[47:32]),
    .b(inputs[15:0]),
    .O0(BIT_ALU_inst0_O0),
    .O1(BIT_ALU_inst0_O1),
    .O2(BIT_ALU_inst0_O2),
    .O3(BIT_ALU_inst0_O3),
    .O4(BIT_ALU_inst0_O4),
    .O5(BIT_ALU_inst0_O5),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
Cond Cond_inst0 (
    .code(inst[6:2]),
    .alu(GTE_inst0_O1),
    .Z(GTE_inst0_O2),
    .N(GTE_inst0_O3),
    .C(GTE_inst0_O4),
    .V(GTE_inst0_O5),
    .O(Cond_inst0_O),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
Cond Cond_inst1 (
    .code(inst[11:7]),
    .alu(LTE_inst0_O1),
    .Z(LTE_inst0_O2),
    .N(LTE_inst0_O3),
    .C(LTE_inst0_O4),
    .V(LTE_inst0_O5),
    .O(Cond_inst1_O),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
Cond Cond_inst2 (
    .code(inst[16:12]),
    .alu(SUB_inst0_O1),
    .Z(SUB_inst0_O2),
    .N(SUB_inst0_O3),
    .C(SUB_inst0_O4),
    .V(SUB_inst0_O5),
    .O(Cond_inst2_O),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
GTE GTE_inst0 (
    .signed_(inst[46]),
    .a(inputs[47:32]),
    .b(inputs[15:0]),
    .O0(GTE_inst0_O0),
    .O1(GTE_inst0_O1),
    .O2(GTE_inst0_O2),
    .O3(GTE_inst0_O3),
    .O4(GTE_inst0_O4),
    .O5(GTE_inst0_O5),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
LTE LTE_inst0 (
    .signed_(inst[47]),
    .a(inputs[47:32]),
    .b(inputs[15:0]),
    .O0(LTE_inst0_O0),
    .O1(LTE_inst0_O1),
    .O2(LTE_inst0_O2),
    .O3(LTE_inst0_O3),
    .O4(LTE_inst0_O4),
    .O5(LTE_inst0_O5),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
LUT LUT_inst0 (
    .lut(inst[56:49]),
    .bit0(inputs[48]),
    .bit1(inputs[49]),
    .bit2(inputs[50]),
    .O(LUT_inst0_O),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
MUL MUL_inst0 (
    .instr(inst[18:17]),
    .signed_(inst[45]),
    .a(inputs[47:32]),
    .b(Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out),
    .O(MUL_inst0_O),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Cond_inst0_O),
    .in1(Cond_inst0_O),
    .sel(magma_Bits_3_eq_inst0_out),
    .out(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst0$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(Cond_inst1_O),
    .sel(magma_Bits_3_eq_inst1_out),
    .out(Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst1$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(Cond_inst2_O),
    .sel(magma_Bits_3_eq_inst2_out),
    .out(Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst2$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(inst[35]),
    .sel(magma_Bits_3_eq_inst3_out),
    .out(Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(1)
) Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join (
    .in0(Mux2xBit_inst3$coreir_commonlib_mux2x1_inst0$_join_out[0]),
    .in1(LUT_inst0_O),
    .sel(magma_Bits_3_eq_inst4_out),
    .out(Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst0_I0_in),
    .in1(Mux2xBits16_inst0_I1_in),
    .sel(magma_Bits_1_eq_inst0_out),
    .out(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
mantle_wire__typeBitIn16 Mux2xBits16_inst0_I0 (
    .in(Mux2xBits16_inst0_I0_in),
    .out(inst[34:19])
);
mantle_wire__typeBitIn16 Mux2xBits16_inst0_I1 (
    .in(Mux2xBits16_inst0_I1_in),
    .out(inst[34:19])
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(Mux2xBits16_inst1_I1_in),
    .sel(magma_Bits_1_eq_inst1_out),
    .out(Mux2xBits16_inst1$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst10$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst9$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(ABSD_inst0_O0),
    .sel(magma_Bits_4_eq_inst6_out),
    .out(Mux2xBits16_inst10$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst11$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst10$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(SHR_inst0_O0),
    .sel(magma_Bits_4_eq_inst7_out),
    .out(Mux2xBits16_inst11$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst12$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst11$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(BIT_ALU_inst0_O0),
    .sel(magma_Bits_4_eq_inst8_out),
    .out(Mux2xBits16_inst12$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst13$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst12$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(ADD_inst1_O0),
    .sel(magma_Bits_4_eq_inst9_out),
    .out(Mux2xBits16_inst13$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst14$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst13$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(MUL_inst0_O),
    .sel(magma_Bits_4_eq_inst10_out),
    .out(Mux2xBits16_inst14$coreir_commonlib_mux2x16_inst0$_join_out)
);
mantle_wire__typeBit16 Mux2xBits16_inst14_O (
    .in(Mux2xBits16_inst14$coreir_commonlib_mux2x16_inst0$_join_out),
    .out(Mux2xBits16_inst14_O_out)
);
mantle_wire__typeBitIn16 Mux2xBits16_inst1_I1 (
    .in(Mux2xBits16_inst1_I1_in),
    .out(inputs[15:0])
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst2_I0_in),
    .in1(Mux2xBits16_inst2_I1_in),
    .sel(magma_Bits_1_eq_inst2_out),
    .out(Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_out)
);
mantle_wire__typeBitIn16 Mux2xBits16_inst2_I0 (
    .in(Mux2xBits16_inst2_I0_in),
    .out(inst[34:19])
);
mantle_wire__typeBitIn16 Mux2xBits16_inst2_I1 (
    .in(Mux2xBits16_inst2_I1_in),
    .out(inst[34:19])
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst2$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(ADD_inst0_O0),
    .sel(magma_Bits_1_eq_inst3_out),
    .out(Mux2xBits16_inst3$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join (
    .in0(ADD_inst0_O0),
    .in1(ADD_inst0_O0),
    .sel(magma_Bits_4_eq_inst0_out),
    .out(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst5$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst4$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(GTE_inst0_O0),
    .sel(magma_Bits_4_eq_inst1_out),
    .out(Mux2xBits16_inst5$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst6$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst5$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(Mux_inst0$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out),
    .sel(magma_Bits_4_eq_inst2_out),
    .out(Mux2xBits16_inst6$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst6$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(LTE_inst0_O0),
    .sel(magma_Bits_4_eq_inst3_out),
    .out(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst8$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst7$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(SUB_inst0_O0),
    .sel(magma_Bits_4_eq_inst4_out),
    .out(Mux2xBits16_inst8$coreir_commonlib_mux2x16_inst0$_join_out)
);
coreir_mux #(
    .width(16)
) Mux2xBits16_inst9$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux2xBits16_inst8$coreir_commonlib_mux2x16_inst0$_join_out),
    .in1(Mux2xBits16_inst9_I1_in),
    .sel(magma_Bits_4_eq_inst5_out),
    .out(Mux2xBits16_inst9$coreir_commonlib_mux2x16_inst0$_join_out)
);
mantle_wire__typeBitIn16 Mux2xBits16_inst9_I1 (
    .in(Mux2xBits16_inst9_I1_in),
    .out(inst[34:19])
);
coreir_mux #(
    .width(16)
) Mux_inst0$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join (
    .in0(Mux_inst0_a_in),
    .in1(Mux_inst0_b_in),
    .sel(inputs[48]),
    .out(Mux_inst0$Mux2xBits16_inst0$coreir_commonlib_mux2x16_inst0$_join_out)
);
mantle_wire__typeBitIn16 Mux_inst0_a (
    .in(Mux_inst0_a_in),
    .out(inputs[31:16])
);
mantle_wire__typeBitIn16 Mux_inst0_b (
    .in(Mux_inst0_b_in),
    .out(inputs[47:32])
);
SHR SHR_inst0 (
    .signed_(inst[48]),
    .a(inputs[47:32]),
    .b(inputs[15:0]),
    .O0(SHR_inst0_O0),
    .O1(SHR_inst0_O1),
    .O2(SHR_inst0_O2),
    .O3(SHR_inst0_O3),
    .O4(SHR_inst0_O4),
    .O5(SHR_inst0_O5),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
SUB SUB_inst0 (
    .a(inputs[31:16]),
    .b(inputs[47:32]),
    .O0(SUB_inst0_O0),
    .O1(SUB_inst0_O1),
    .O2(SUB_inst0_O2),
    .O3(SUB_inst0_O3),
    .O4(SUB_inst0_O4),
    .O5(SUB_inst0_O5),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
coreir_const #(
    .value(1'h0),
    .width(1)
) const_0_1 (
    .out(const_0_1_out)
);
coreir_const #(
    .value(3'h0),
    .width(3)
) const_0_3 (
    .out(const_0_3_out)
);
coreir_const #(
    .value(4'h0),
    .width(4)
) const_0_4 (
    .out(const_0_4_out)
);
coreir_const #(
    .value(4'ha),
    .width(4)
) const_10_4 (
    .out(const_10_4_out)
);
coreir_const #(
    .value(1'h1),
    .width(1)
) const_1_1 (
    .out(const_1_1_out)
);
coreir_const #(
    .value(3'h1),
    .width(3)
) const_1_3 (
    .out(const_1_3_out)
);
coreir_const #(
    .value(4'h1),
    .width(4)
) const_1_4 (
    .out(const_1_4_out)
);
coreir_const #(
    .value(3'h2),
    .width(3)
) const_2_3 (
    .out(const_2_3_out)
);
coreir_const #(
    .value(4'h2),
    .width(4)
) const_2_4 (
    .out(const_2_4_out)
);
coreir_const #(
    .value(3'h3),
    .width(3)
) const_3_3 (
    .out(const_3_3_out)
);
coreir_const #(
    .value(4'h3),
    .width(4)
) const_3_4 (
    .out(const_3_4_out)
);
coreir_const #(
    .value(3'h4),
    .width(3)
) const_4_3 (
    .out(const_4_3_out)
);
coreir_const #(
    .value(4'h4),
    .width(4)
) const_4_4 (
    .out(const_4_4_out)
);
coreir_const #(
    .value(4'h5),
    .width(4)
) const_5_4 (
    .out(const_5_4_out)
);
coreir_const #(
    .value(4'h6),
    .width(4)
) const_6_4 (
    .out(const_6_4_out)
);
coreir_const #(
    .value(4'h7),
    .width(4)
) const_7_4 (
    .out(const_7_4_out)
);
coreir_const #(
    .value(4'h8),
    .width(4)
) const_8_4 (
    .out(const_8_4_out)
);
coreir_const #(
    .value(4'h9),
    .width(4)
) const_9_4 (
    .out(const_9_4_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst0 (
    .in0(inst[36]),
    .in1(const_0_1_out),
    .out(magma_Bits_1_eq_inst0_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst1 (
    .in0(inst[36]),
    .in1(const_1_1_out),
    .out(magma_Bits_1_eq_inst1_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst2 (
    .in0(inst[37]),
    .in1(const_0_1_out),
    .out(magma_Bits_1_eq_inst2_out)
);
coreir_eq #(
    .width(1)
) magma_Bits_1_eq_inst3 (
    .in0(inst[37]),
    .in1(const_1_1_out),
    .out(magma_Bits_1_eq_inst3_out)
);
coreir_eq #(
    .width(3)
) magma_Bits_3_eq_inst0 (
    .in0(inst[44:42]),
    .in1(const_0_3_out),
    .out(magma_Bits_3_eq_inst0_out)
);
coreir_eq #(
    .width(3)
) magma_Bits_3_eq_inst1 (
    .in0(inst[44:42]),
    .in1(const_1_3_out),
    .out(magma_Bits_3_eq_inst1_out)
);
coreir_eq #(
    .width(3)
) magma_Bits_3_eq_inst2 (
    .in0(inst[44:42]),
    .in1(const_2_3_out),
    .out(magma_Bits_3_eq_inst2_out)
);
coreir_eq #(
    .width(3)
) magma_Bits_3_eq_inst3 (
    .in0(inst[44:42]),
    .in1(const_3_3_out),
    .out(magma_Bits_3_eq_inst3_out)
);
coreir_eq #(
    .width(3)
) magma_Bits_3_eq_inst4 (
    .in0(inst[44:42]),
    .in1(const_4_3_out),
    .out(magma_Bits_3_eq_inst4_out)
);
coreir_eq #(
    .width(4)
) magma_Bits_4_eq_inst0 (
    .in0(inst[41:38]),
    .in1(const_0_4_out),
    .out(magma_Bits_4_eq_inst0_out)
);
coreir_eq #(
    .width(4)
) magma_Bits_4_eq_inst1 (
    .in0(inst[41:38]),
    .in1(const_1_4_out),
    .out(magma_Bits_4_eq_inst1_out)
);
coreir_eq #(
    .width(4)
) magma_Bits_4_eq_inst10 (
    .in0(inst[41:38]),
    .in1(const_10_4_out),
    .out(magma_Bits_4_eq_inst10_out)
);
coreir_eq #(
    .width(4)
) magma_Bits_4_eq_inst2 (
    .in0(inst[41:38]),
    .in1(const_2_4_out),
    .out(magma_Bits_4_eq_inst2_out)
);
coreir_eq #(
    .width(4)
) magma_Bits_4_eq_inst3 (
    .in0(inst[41:38]),
    .in1(const_3_4_out),
    .out(magma_Bits_4_eq_inst3_out)
);
coreir_eq #(
    .width(4)
) magma_Bits_4_eq_inst4 (
    .in0(inst[41:38]),
    .in1(const_4_4_out),
    .out(magma_Bits_4_eq_inst4_out)
);
coreir_eq #(
    .width(4)
) magma_Bits_4_eq_inst5 (
    .in0(inst[41:38]),
    .in1(const_5_4_out),
    .out(magma_Bits_4_eq_inst5_out)
);
coreir_eq #(
    .width(4)
) magma_Bits_4_eq_inst6 (
    .in0(inst[41:38]),
    .in1(const_6_4_out),
    .out(magma_Bits_4_eq_inst6_out)
);
coreir_eq #(
    .width(4)
) magma_Bits_4_eq_inst7 (
    .in0(inst[41:38]),
    .in1(const_7_4_out),
    .out(magma_Bits_4_eq_inst7_out)
);
coreir_eq #(
    .width(4)
) magma_Bits_4_eq_inst8 (
    .in0(inst[41:38]),
    .in1(const_8_4_out),
    .out(magma_Bits_4_eq_inst8_out)
);
coreir_eq #(
    .width(4)
) magma_Bits_4_eq_inst9 (
    .in0(inst[41:38]),
    .in1(const_9_4_out),
    .out(magma_Bits_4_eq_inst9_out)
);
assign O = {Mux2xBit_inst4$coreir_commonlib_mux2x1_inst0$_join_out[0],Mux2xBits16_inst14_O_out[15:0]};
endmodule

module WrappedPE (
    input [56:0] inst,
    input [15:0] inputs0,
    input [15:0] inputs1,
    input [15:0] inputs2,
    input inputs3,
    input inputs4,
    input inputs5,
    input clk_en,
    output [15:0] O0,
    output O1,
    input CLK,
    input ASYNCRESET
);
wire [16:0] PE_inst0$PE_gen_inst0_O;
wire [15:0] PE_inst0$self_O0_in;
wire [15:0] PE_inst0$self_inputs0_out;
wire [15:0] PE_inst0$self_inputs1_out;
wire [15:0] PE_inst0$self_inputs2_out;
wire [50:0] PE_inst0$PE_gen_inst0_inputs;
assign PE_inst0$PE_gen_inst0_inputs = {inputs5,inputs4,inputs3,PE_inst0$self_inputs2_out[15:0],PE_inst0$self_inputs1_out[15:0],PE_inst0$self_inputs0_out[15:0]};
PE_gen PE_inst0$PE_gen_inst0 (
    .inst(inst),
    .inputs(PE_inst0$PE_gen_inst0_inputs),
    .clk_en(clk_en),
    .O(PE_inst0$PE_gen_inst0_O),
    .CLK(CLK),
    .ASYNCRESET(ASYNCRESET)
);
mantle_wire__typeBitIn16 PE_inst0$self_O0 (
    .in(PE_inst0$self_O0_in),
    .out(PE_inst0$PE_gen_inst0_O[15:0])
);
mantle_wire__typeBit16 PE_inst0$self_inputs0 (
    .in(inputs0),
    .out(PE_inst0$self_inputs0_out)
);
mantle_wire__typeBit16 PE_inst0$self_inputs1 (
    .in(inputs1),
    .out(PE_inst0$self_inputs1_out)
);
mantle_wire__typeBit16 PE_inst0$self_inputs2 (
    .in(inputs2),
    .out(PE_inst0$self_inputs2_out)
);
assign O0 = PE_inst0$self_O0_in;
assign O1 = PE_inst0$PE_gen_inst0_O[16];
endmodule

module PE_unq1 (
    input clk,
    input [7:0] config_config_addr,
    input [31:0] config_config_data,
    input [0:0] config_read,
    input [0:0] config_write,
    input [15:0] inputs0,
    input [15:0] inputs1,
    input [15:0] inputs2,
    input [0:0] inputs3,
    input [0:0] inputs4,
    input [0:0] inputs5,
    output [15:0] pe_outputs_0,
    output [0:0] pe_outputs_1,
    output [31:0] read_config_data,
    input reset,
    input [0:0] stall
);
wire [0:0] Invert1_inst0_out;
wire [31:0] MuxWrapper_2_32_inst0$Mux2x32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
wire [15:0] WrappedPE_inst0_O0;
wire WrappedPE_inst0_O1;
wire [31:0] config_reg_0_O;
wire [31:0] config_reg_1_O;
wire [31:0] inst_0_inst0_O;
wire [31:0] inst_1_inst0_O;
coreir_not #(
    .width(1)
) Invert1_inst0 (
    .in(stall),
    .out(Invert1_inst0_out)
);
coreir_mux #(
    .width(32)
) MuxWrapper_2_32_inst0$Mux2x32_inst0$coreir_commonlib_mux2x32_inst0$_join (
    .in0(config_reg_0_O),
    .in1(config_reg_1_O),
    .sel(config_config_addr[0]),
    .out(MuxWrapper_2_32_inst0$Mux2x32_inst0$coreir_commonlib_mux2x32_inst0$_join_out)
);
wire [56:0] WrappedPE_inst0_inst;
assign WrappedPE_inst0_inst = {inst_1_inst0_O[24:0],inst_0_inst0_O[31:0]};
WrappedPE WrappedPE_inst0 (
    .inst(WrappedPE_inst0_inst),
    .inputs0(inputs0),
    .inputs1(inputs1),
    .inputs2(inputs2),
    .inputs3(inputs3[0]),
    .inputs4(inputs4[0]),
    .inputs5(inputs5[0]),
    .clk_en(Invert1_inst0_out[0]),
    .O0(WrappedPE_inst0_O0),
    .O1(WrappedPE_inst0_O1),
    .CLK(clk),
    .ASYNCRESET(reset)
);
ConfigRegister_32_8_32_0 config_reg_0 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_0_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
ConfigRegister_32_8_32_1 config_reg_1 (
    .clk(clk),
    .reset(reset),
    .O(config_reg_1_O),
    .config_addr(config_config_addr),
    .config_data(config_config_data),
    .config_en(config_write[0])
);
inst_0 inst_0_inst0 (
    .I(config_reg_0_O),
    .O(inst_0_inst0_O)
);
inst_1 inst_1_inst0 (
    .I(config_reg_1_O),
    .O(inst_1_inst0_O)
);
assign pe_outputs_0 = WrappedPE_inst0_O0;
assign pe_outputs_1 = WrappedPE_inst0_O1;
assign read_config_data = MuxWrapper_2_32_inst0$Mux2x32_inst0$coreir_commonlib_mux2x32_inst0$_join_out;
endmodule

module Tile_PE (
    input [0:0] SB_T0_EAST_SB_IN_B1,
    input [15:0] SB_T0_EAST_SB_IN_B16,
    output [0:0] SB_T0_EAST_SB_OUT_B1,
    output [15:0] SB_T0_EAST_SB_OUT_B16,
    input [0:0] SB_T0_NORTH_SB_IN_B1,
    input [15:0] SB_T0_NORTH_SB_IN_B16,
    output [0:0] SB_T0_NORTH_SB_OUT_B1,
    output [15:0] SB_T0_NORTH_SB_OUT_B16,
    input [0:0] SB_T0_SOUTH_SB_IN_B1,
    input [15:0] SB_T0_SOUTH_SB_IN_B16,
    output [0:0] SB_T0_SOUTH_SB_OUT_B1,
    output [15:0] SB_T0_SOUTH_SB_OUT_B16,
    input [0:0] SB_T0_WEST_SB_IN_B1,
    input [15:0] SB_T0_WEST_SB_IN_B16,
    output [0:0] SB_T0_WEST_SB_OUT_B1,
    output [15:0] SB_T0_WEST_SB_OUT_B16,
    input [0:0] SB_T1_EAST_SB_IN_B1,
    input [15:0] SB_T1_EAST_SB_IN_B16,
    output [0:0] SB_T1_EAST_SB_OUT_B1,
    output [15:0] SB_T1_EAST_SB_OUT_B16,
    input [0:0] SB_T1_NORTH_SB_IN_B1,
    input [15:0] SB_T1_NORTH_SB_IN_B16,
    output [0:0] SB_T1_NORTH_SB_OUT_B1,
    output [15:0] SB_T1_NORTH_SB_OUT_B16,
    input [0:0] SB_T1_SOUTH_SB_IN_B1,
    input [15:0] SB_T1_SOUTH_SB_IN_B16,
    output [0:0] SB_T1_SOUTH_SB_OUT_B1,
    output [15:0] SB_T1_SOUTH_SB_OUT_B16,
    input [0:0] SB_T1_WEST_SB_IN_B1,
    input [15:0] SB_T1_WEST_SB_IN_B16,
    output [0:0] SB_T1_WEST_SB_OUT_B1,
    output [15:0] SB_T1_WEST_SB_OUT_B16,
    input [0:0] SB_T2_EAST_SB_IN_B1,
    input [15:0] SB_T2_EAST_SB_IN_B16,
    output [0:0] SB_T2_EAST_SB_OUT_B1,
    output [15:0] SB_T2_EAST_SB_OUT_B16,
    input [0:0] SB_T2_NORTH_SB_IN_B1,
    input [15:0] SB_T2_NORTH_SB_IN_B16,
    output [0:0] SB_T2_NORTH_SB_OUT_B1,
    output [15:0] SB_T2_NORTH_SB_OUT_B16,
    input [0:0] SB_T2_SOUTH_SB_IN_B1,
    input [15:0] SB_T2_SOUTH_SB_IN_B16,
    output [0:0] SB_T2_SOUTH_SB_OUT_B1,
    output [15:0] SB_T2_SOUTH_SB_OUT_B16,
    input [0:0] SB_T2_WEST_SB_IN_B1,
    input [15:0] SB_T2_WEST_SB_IN_B16,
    output [0:0] SB_T2_WEST_SB_OUT_B1,
    output [15:0] SB_T2_WEST_SB_OUT_B16,
    input [0:0] SB_T3_EAST_SB_IN_B1,
    input [15:0] SB_T3_EAST_SB_IN_B16,
    output [0:0] SB_T3_EAST_SB_OUT_B1,
    output [15:0] SB_T3_EAST_SB_OUT_B16,
    input [0:0] SB_T3_NORTH_SB_IN_B1,
    input [15:0] SB_T3_NORTH_SB_IN_B16,
    output [0:0] SB_T3_NORTH_SB_OUT_B1,
    output [15:0] SB_T3_NORTH_SB_OUT_B16,
    input [0:0] SB_T3_SOUTH_SB_IN_B1,
    input [15:0] SB_T3_SOUTH_SB_IN_B16,
    output [0:0] SB_T3_SOUTH_SB_OUT_B1,
    output [15:0] SB_T3_SOUTH_SB_OUT_B16,
    input [0:0] SB_T3_WEST_SB_IN_B1,
    input [15:0] SB_T3_WEST_SB_IN_B16,
    output [0:0] SB_T3_WEST_SB_OUT_B1,
    output [15:0] SB_T3_WEST_SB_OUT_B16,
    input [0:0] SB_T4_EAST_SB_IN_B1,
    input [15:0] SB_T4_EAST_SB_IN_B16,
    output [0:0] SB_T4_EAST_SB_OUT_B1,
    output [15:0] SB_T4_EAST_SB_OUT_B16,
    input [0:0] SB_T4_NORTH_SB_IN_B1,
    input [15:0] SB_T4_NORTH_SB_IN_B16,
    output [0:0] SB_T4_NORTH_SB_OUT_B1,
    output [15:0] SB_T4_NORTH_SB_OUT_B16,
    input [0:0] SB_T4_SOUTH_SB_IN_B1,
    input [15:0] SB_T4_SOUTH_SB_IN_B16,
    output [0:0] SB_T4_SOUTH_SB_OUT_B1,
    output [15:0] SB_T4_SOUTH_SB_OUT_B16,
    input [0:0] SB_T4_WEST_SB_IN_B1,
    input [15:0] SB_T4_WEST_SB_IN_B16,
    output [0:0] SB_T4_WEST_SB_OUT_B1,
    output [15:0] SB_T4_WEST_SB_OUT_B16,
    input clk,
    output clk_out,
    input clk_pass_through,
    output clk_pass_through_out_bot,
    output clk_pass_through_out_right,
    input [31:0] config_config_addr,
    input [31:0] config_config_data,
    output [31:0] config_out_config_addr,
    output [31:0] config_out_config_data,
    output [0:0] config_out_read,
    output [0:0] config_out_write,
    input [0:0] config_read,
    input [0:0] config_write,
    output [8:0] hi,
    output [7:0] lo,
    output [31:0] read_config_data,
    input [31:0] read_config_data_in,
    input reset,
    output reset_out,
    input [0:0] stall,
    output [0:0] stall_out,
    input [15:0] tile_id
);
wire [15:0] CB_inputs0_O;
wire [31:0] CB_inputs0_read_config_data;
wire [7:0] CB_inputs0_config_config_addr_in;
wire [15:0] CB_inputs1_O;
wire [31:0] CB_inputs1_read_config_data;
wire [7:0] CB_inputs1_config_config_addr_in;
wire [15:0] CB_inputs2_O;
wire [31:0] CB_inputs2_read_config_data;
wire [7:0] CB_inputs2_config_config_addr_in;
wire [0:0] CB_inputs3_O;
wire [31:0] CB_inputs3_read_config_data;
wire [7:0] CB_inputs3_config_config_addr_in;
wire [0:0] CB_inputs4_O;
wire [31:0] CB_inputs4_read_config_data;
wire [7:0] CB_inputs4_config_config_addr_in;
wire [0:0] CB_inputs5_O;
wire [31:0] CB_inputs5_read_config_data;
wire [7:0] CB_inputs5_config_config_addr_in;
wire DECODE_FEATURE_0_O;
wire DECODE_FEATURE_1_O;
wire DECODE_FEATURE_2_O;
wire DECODE_FEATURE_3_O;
wire DECODE_FEATURE_4_O;
wire DECODE_FEATURE_5_O;
wire DECODE_FEATURE_6_O;
wire DECODE_FEATURE_7_O;
wire DECODE_FEATURE_8_O;
wire FEATURE_AND_0_out;
wire FEATURE_AND_1_out;
wire FEATURE_AND_2_out;
wire FEATURE_AND_3_out;
wire FEATURE_AND_4_out;
wire FEATURE_AND_5_out;
wire FEATURE_AND_6_out;
wire FEATURE_AND_7_out;
wire FEATURE_AND_8_out;
wire [15:0] PE_inst0_pe_outputs_0;
wire [0:0] PE_inst0_pe_outputs_1;
wire [31:0] PE_inst0_read_config_data;
wire [7:0] PE_inst0_config_config_addr_in;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T0_EAST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T0_NORTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T0_SOUTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T0_WEST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T1_EAST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T1_NORTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T1_SOUTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T1_WEST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T2_EAST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T2_NORTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T2_SOUTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T2_WEST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T3_EAST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T3_NORTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T3_SOUTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T3_WEST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T4_EAST_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T4_NORTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T4_SOUTH_SB_OUT_B16;
wire [15:0] SB_ID0_5TRACKS_B16_PE_SB_T4_WEST_SB_OUT_B16;
wire [31:0] SB_ID0_5TRACKS_B16_PE_read_config_data;
wire [7:0] SB_ID0_5TRACKS_B16_PE_config_config_addr_in;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_OUT_B1;
wire [0:0] SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_OUT_B1;
wire [31:0] SB_ID0_5TRACKS_B1_PE_read_config_data;
wire [7:0] SB_ID0_5TRACKS_B1_PE_config_config_addr_in;
wire [0:0] WIRE_SB_T0_EAST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T0_EAST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T0_NORTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T0_NORTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T0_SOUTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T0_SOUTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T0_WEST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T0_WEST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T1_EAST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T1_EAST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T1_NORTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T1_NORTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T1_SOUTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T1_SOUTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T1_WEST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T1_WEST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T2_EAST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T2_EAST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T2_NORTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T2_NORTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T2_SOUTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T2_SOUTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T2_WEST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T2_WEST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T3_EAST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T3_EAST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T3_NORTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T3_NORTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T3_SOUTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T3_SOUTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T3_WEST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T3_WEST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T4_EAST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T4_EAST_SB_IN_B16_O;
wire [0:0] WIRE_SB_T4_NORTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T4_NORTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T4_SOUTH_SB_IN_B1_O;
wire [15:0] WIRE_SB_T4_SOUTH_SB_IN_B16_O;
wire [0:0] WIRE_SB_T4_WEST_SB_IN_B1_O;
wire [15:0] WIRE_SB_T4_WEST_SB_IN_B16_O;
wire and_inst0_out;
wire and_inst1_out;
wire [7:0] const_0_8_out;
wire [8:0] const_511_9_out;
wire coreir_eq_16_inst0_out;
wire [31:0] read_config_data_or_inst0_out;
wire [31:0] read_data_mux_O;
wire [7:0] read_data_mux_S_in;
wire [31:0] self_config_config_addr_out;
CB_inputs0 CB_inputs0 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .O(CB_inputs0_O),
    .clk(clk),
    .config_config_addr(CB_inputs0_config_config_addr_in),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_1_out),
    .read_config_data(CB_inputs0_read_config_data),
    .reset(reset)
);
mantle_wire__typeBitIn8 CB_inputs0_config_config_addr (
    .in(CB_inputs0_config_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
CB_inputs1 CB_inputs1 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .O(CB_inputs1_O),
    .clk(clk),
    .config_config_addr(CB_inputs1_config_config_addr_in),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_2_out),
    .read_config_data(CB_inputs1_read_config_data),
    .reset(reset)
);
mantle_wire__typeBitIn8 CB_inputs1_config_config_addr (
    .in(CB_inputs1_config_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
CB_inputs2 CB_inputs2 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B16_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B16_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B16_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B16_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B16_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B16_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B16_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B16_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B16_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B16_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B16_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B16_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B16_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B16_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B16_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B16_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B16_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B16_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B16_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B16_O),
    .O(CB_inputs2_O),
    .clk(clk),
    .config_config_addr(CB_inputs2_config_config_addr_in),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_3_out),
    .read_config_data(CB_inputs2_read_config_data),
    .reset(reset)
);
mantle_wire__typeBitIn8 CB_inputs2_config_config_addr (
    .in(CB_inputs2_config_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
CB_inputs3 CB_inputs3 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .O(CB_inputs3_O),
    .clk(clk),
    .config_config_addr(CB_inputs3_config_config_addr_in),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_4_out),
    .read_config_data(CB_inputs3_read_config_data),
    .reset(reset)
);
mantle_wire__typeBitIn8 CB_inputs3_config_config_addr (
    .in(CB_inputs3_config_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
CB_inputs4 CB_inputs4 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .O(CB_inputs4_O),
    .clk(clk),
    .config_config_addr(CB_inputs4_config_config_addr_in),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_5_out),
    .read_config_data(CB_inputs4_read_config_data),
    .reset(reset)
);
mantle_wire__typeBitIn8 CB_inputs4_config_config_addr (
    .in(CB_inputs4_config_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
CB_inputs5 CB_inputs5 (
    .I_0(WIRE_SB_T0_NORTH_SB_IN_B1_O),
    .I_1(WIRE_SB_T0_SOUTH_SB_IN_B1_O),
    .I_10(WIRE_SB_T2_EAST_SB_IN_B1_O),
    .I_11(WIRE_SB_T2_WEST_SB_IN_B1_O),
    .I_12(WIRE_SB_T3_NORTH_SB_IN_B1_O),
    .I_13(WIRE_SB_T3_SOUTH_SB_IN_B1_O),
    .I_14(WIRE_SB_T3_EAST_SB_IN_B1_O),
    .I_15(WIRE_SB_T3_WEST_SB_IN_B1_O),
    .I_16(WIRE_SB_T4_NORTH_SB_IN_B1_O),
    .I_17(WIRE_SB_T4_SOUTH_SB_IN_B1_O),
    .I_18(WIRE_SB_T4_EAST_SB_IN_B1_O),
    .I_19(WIRE_SB_T4_WEST_SB_IN_B1_O),
    .I_2(WIRE_SB_T0_EAST_SB_IN_B1_O),
    .I_3(WIRE_SB_T0_WEST_SB_IN_B1_O),
    .I_4(WIRE_SB_T1_NORTH_SB_IN_B1_O),
    .I_5(WIRE_SB_T1_SOUTH_SB_IN_B1_O),
    .I_6(WIRE_SB_T1_EAST_SB_IN_B1_O),
    .I_7(WIRE_SB_T1_WEST_SB_IN_B1_O),
    .I_8(WIRE_SB_T2_NORTH_SB_IN_B1_O),
    .I_9(WIRE_SB_T2_SOUTH_SB_IN_B1_O),
    .O(CB_inputs5_O),
    .clk(clk),
    .config_config_addr(CB_inputs5_config_config_addr_in),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_6_out),
    .read_config_data(CB_inputs5_read_config_data),
    .reset(reset)
);
mantle_wire__typeBitIn8 CB_inputs5_config_config_addr (
    .in(CB_inputs5_config_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
Decode08 DECODE_FEATURE_0 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_0_O)
);
Decode18 DECODE_FEATURE_1 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_1_O)
);
Decode28 DECODE_FEATURE_2 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_2_O)
);
Decode38 DECODE_FEATURE_3 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_3_O)
);
Decode48 DECODE_FEATURE_4 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_4_O)
);
Decode58 DECODE_FEATURE_5 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_5_O)
);
Decode68 DECODE_FEATURE_6 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_6_O)
);
Decode78 DECODE_FEATURE_7 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_7_O)
);
Decode88 DECODE_FEATURE_8 (
    .I(self_config_config_addr_out[23:16]),
    .O(DECODE_FEATURE_8_O)
);
corebit_and FEATURE_AND_0 (
    .in0(DECODE_FEATURE_0_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_0_out)
);
corebit_and FEATURE_AND_1 (
    .in0(DECODE_FEATURE_1_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_1_out)
);
corebit_and FEATURE_AND_2 (
    .in0(DECODE_FEATURE_2_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_2_out)
);
corebit_and FEATURE_AND_3 (
    .in0(DECODE_FEATURE_3_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_3_out)
);
corebit_and FEATURE_AND_4 (
    .in0(DECODE_FEATURE_4_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_4_out)
);
corebit_and FEATURE_AND_5 (
    .in0(DECODE_FEATURE_5_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_5_out)
);
corebit_and FEATURE_AND_6 (
    .in0(DECODE_FEATURE_6_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_6_out)
);
corebit_and FEATURE_AND_7 (
    .in0(DECODE_FEATURE_7_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_7_out)
);
corebit_and FEATURE_AND_8 (
    .in0(DECODE_FEATURE_8_O),
    .in1(and_inst1_out),
    .out(FEATURE_AND_8_out)
);
PE_unq1 PE_inst0 (
    .clk(clk),
    .config_config_addr(PE_inst0_config_config_addr_in),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_0_out),
    .inputs0(CB_inputs0_O),
    .inputs1(CB_inputs1_O),
    .inputs2(CB_inputs2_O),
    .inputs3(CB_inputs3_O),
    .inputs4(CB_inputs4_O),
    .inputs5(CB_inputs5_O),
    .pe_outputs_0(PE_inst0_pe_outputs_0),
    .pe_outputs_1(PE_inst0_pe_outputs_1),
    .read_config_data(PE_inst0_read_config_data),
    .reset(reset),
    .stall(stall)
);
mantle_wire__typeBitIn8 PE_inst0_config_config_addr (
    .in(PE_inst0_config_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
SB_ID0_5TRACKS_B16_PE SB_ID0_5TRACKS_B16_PE (
    .SB_T0_EAST_SB_IN_B16(SB_T0_EAST_SB_IN_B16),
    .SB_T0_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B16(SB_T0_NORTH_SB_IN_B16),
    .SB_T0_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B16(SB_T0_SOUTH_SB_IN_B16),
    .SB_T0_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B16(SB_T0_WEST_SB_IN_B16),
    .SB_T0_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B16(SB_T1_EAST_SB_IN_B16),
    .SB_T1_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B16(SB_T1_NORTH_SB_IN_B16),
    .SB_T1_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B16(SB_T1_SOUTH_SB_IN_B16),
    .SB_T1_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B16(SB_T1_WEST_SB_IN_B16),
    .SB_T1_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B16(SB_T2_EAST_SB_IN_B16),
    .SB_T2_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B16(SB_T2_NORTH_SB_IN_B16),
    .SB_T2_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B16(SB_T2_SOUTH_SB_IN_B16),
    .SB_T2_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B16(SB_T2_WEST_SB_IN_B16),
    .SB_T2_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B16(SB_T3_EAST_SB_IN_B16),
    .SB_T3_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B16(SB_T3_NORTH_SB_IN_B16),
    .SB_T3_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B16(SB_T3_SOUTH_SB_IN_B16),
    .SB_T3_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B16(SB_T3_WEST_SB_IN_B16),
    .SB_T3_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B16(SB_T4_EAST_SB_IN_B16),
    .SB_T4_EAST_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B16(SB_T4_NORTH_SB_IN_B16),
    .SB_T4_NORTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B16(SB_T4_SOUTH_SB_IN_B16),
    .SB_T4_SOUTH_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B16(SB_T4_WEST_SB_IN_B16),
    .SB_T4_WEST_SB_OUT_B16(SB_ID0_5TRACKS_B16_PE_SB_T4_WEST_SB_OUT_B16),
    .clk(clk),
    .config_config_addr(SB_ID0_5TRACKS_B16_PE_config_config_addr_in),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_8_out),
    .pe_outputs_0(PE_inst0_pe_outputs_0),
    .read_config_data(SB_ID0_5TRACKS_B16_PE_read_config_data),
    .reset(reset),
    .stall(stall)
);
mantle_wire__typeBitIn8 SB_ID0_5TRACKS_B16_PE_config_config_addr (
    .in(SB_ID0_5TRACKS_B16_PE_config_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
SB_ID0_5TRACKS_B1_PE SB_ID0_5TRACKS_B1_PE (
    .SB_T0_EAST_SB_IN_B1(SB_T0_EAST_SB_IN_B1),
    .SB_T0_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B1(SB_T0_NORTH_SB_IN_B1),
    .SB_T0_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B1(SB_T0_SOUTH_SB_IN_B1),
    .SB_T0_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B1(SB_T0_WEST_SB_IN_B1),
    .SB_T0_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B1(SB_T1_EAST_SB_IN_B1),
    .SB_T1_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B1(SB_T1_NORTH_SB_IN_B1),
    .SB_T1_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B1(SB_T1_SOUTH_SB_IN_B1),
    .SB_T1_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B1(SB_T1_WEST_SB_IN_B1),
    .SB_T1_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B1(SB_T2_EAST_SB_IN_B1),
    .SB_T2_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B1(SB_T2_NORTH_SB_IN_B1),
    .SB_T2_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B1(SB_T2_SOUTH_SB_IN_B1),
    .SB_T2_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B1(SB_T2_WEST_SB_IN_B1),
    .SB_T2_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B1(SB_T3_EAST_SB_IN_B1),
    .SB_T3_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B1(SB_T3_NORTH_SB_IN_B1),
    .SB_T3_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B1(SB_T3_SOUTH_SB_IN_B1),
    .SB_T3_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B1(SB_T3_WEST_SB_IN_B1),
    .SB_T3_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B1(SB_T4_EAST_SB_IN_B1),
    .SB_T4_EAST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B1(SB_T4_NORTH_SB_IN_B1),
    .SB_T4_NORTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B1(SB_T4_SOUTH_SB_IN_B1),
    .SB_T4_SOUTH_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B1(SB_T4_WEST_SB_IN_B1),
    .SB_T4_WEST_SB_OUT_B1(SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_OUT_B1),
    .clk(clk),
    .config_config_addr(SB_ID0_5TRACKS_B1_PE_config_config_addr_in),
    .config_config_data(config_config_data),
    .config_read(config_read),
    .config_write(FEATURE_AND_7_out),
    .pe_outputs_1(PE_inst0_pe_outputs_1),
    .read_config_data(SB_ID0_5TRACKS_B1_PE_read_config_data),
    .reset(reset),
    .stall(stall)
);
mantle_wire__typeBitIn8 SB_ID0_5TRACKS_B1_PE_config_config_addr (
    .in(SB_ID0_5TRACKS_B1_PE_config_config_addr_in),
    .out(self_config_config_addr_out[31:24])
);
MuxWrapper_1_1 WIRE_SB_T0_EAST_SB_IN_B1 (
    .I(SB_T0_EAST_SB_IN_B1),
    .O(WIRE_SB_T0_EAST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T0_EAST_SB_IN_B16 (
    .I(SB_T0_EAST_SB_IN_B16),
    .O(WIRE_SB_T0_EAST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T0_NORTH_SB_IN_B1 (
    .I(SB_T0_NORTH_SB_IN_B1),
    .O(WIRE_SB_T0_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T0_NORTH_SB_IN_B16 (
    .I(SB_T0_NORTH_SB_IN_B16),
    .O(WIRE_SB_T0_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T0_SOUTH_SB_IN_B1 (
    .I(SB_T0_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T0_SOUTH_SB_IN_B16 (
    .I(SB_T0_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T0_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T0_WEST_SB_IN_B1 (
    .I(SB_T0_WEST_SB_IN_B1),
    .O(WIRE_SB_T0_WEST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T0_WEST_SB_IN_B16 (
    .I(SB_T0_WEST_SB_IN_B16),
    .O(WIRE_SB_T0_WEST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T1_EAST_SB_IN_B1 (
    .I(SB_T1_EAST_SB_IN_B1),
    .O(WIRE_SB_T1_EAST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T1_EAST_SB_IN_B16 (
    .I(SB_T1_EAST_SB_IN_B16),
    .O(WIRE_SB_T1_EAST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T1_NORTH_SB_IN_B1 (
    .I(SB_T1_NORTH_SB_IN_B1),
    .O(WIRE_SB_T1_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T1_NORTH_SB_IN_B16 (
    .I(SB_T1_NORTH_SB_IN_B16),
    .O(WIRE_SB_T1_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T1_SOUTH_SB_IN_B1 (
    .I(SB_T1_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T1_SOUTH_SB_IN_B16 (
    .I(SB_T1_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T1_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T1_WEST_SB_IN_B1 (
    .I(SB_T1_WEST_SB_IN_B1),
    .O(WIRE_SB_T1_WEST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T1_WEST_SB_IN_B16 (
    .I(SB_T1_WEST_SB_IN_B16),
    .O(WIRE_SB_T1_WEST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T2_EAST_SB_IN_B1 (
    .I(SB_T2_EAST_SB_IN_B1),
    .O(WIRE_SB_T2_EAST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T2_EAST_SB_IN_B16 (
    .I(SB_T2_EAST_SB_IN_B16),
    .O(WIRE_SB_T2_EAST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T2_NORTH_SB_IN_B1 (
    .I(SB_T2_NORTH_SB_IN_B1),
    .O(WIRE_SB_T2_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T2_NORTH_SB_IN_B16 (
    .I(SB_T2_NORTH_SB_IN_B16),
    .O(WIRE_SB_T2_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T2_SOUTH_SB_IN_B1 (
    .I(SB_T2_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T2_SOUTH_SB_IN_B16 (
    .I(SB_T2_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T2_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T2_WEST_SB_IN_B1 (
    .I(SB_T2_WEST_SB_IN_B1),
    .O(WIRE_SB_T2_WEST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T2_WEST_SB_IN_B16 (
    .I(SB_T2_WEST_SB_IN_B16),
    .O(WIRE_SB_T2_WEST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T3_EAST_SB_IN_B1 (
    .I(SB_T3_EAST_SB_IN_B1),
    .O(WIRE_SB_T3_EAST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T3_EAST_SB_IN_B16 (
    .I(SB_T3_EAST_SB_IN_B16),
    .O(WIRE_SB_T3_EAST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T3_NORTH_SB_IN_B1 (
    .I(SB_T3_NORTH_SB_IN_B1),
    .O(WIRE_SB_T3_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T3_NORTH_SB_IN_B16 (
    .I(SB_T3_NORTH_SB_IN_B16),
    .O(WIRE_SB_T3_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T3_SOUTH_SB_IN_B1 (
    .I(SB_T3_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T3_SOUTH_SB_IN_B16 (
    .I(SB_T3_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T3_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T3_WEST_SB_IN_B1 (
    .I(SB_T3_WEST_SB_IN_B1),
    .O(WIRE_SB_T3_WEST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T3_WEST_SB_IN_B16 (
    .I(SB_T3_WEST_SB_IN_B16),
    .O(WIRE_SB_T3_WEST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T4_EAST_SB_IN_B1 (
    .I(SB_T4_EAST_SB_IN_B1),
    .O(WIRE_SB_T4_EAST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T4_EAST_SB_IN_B16 (
    .I(SB_T4_EAST_SB_IN_B16),
    .O(WIRE_SB_T4_EAST_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T4_NORTH_SB_IN_B1 (
    .I(SB_T4_NORTH_SB_IN_B1),
    .O(WIRE_SB_T4_NORTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T4_NORTH_SB_IN_B16 (
    .I(SB_T4_NORTH_SB_IN_B16),
    .O(WIRE_SB_T4_NORTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T4_SOUTH_SB_IN_B1 (
    .I(SB_T4_SOUTH_SB_IN_B1),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T4_SOUTH_SB_IN_B16 (
    .I(SB_T4_SOUTH_SB_IN_B16),
    .O(WIRE_SB_T4_SOUTH_SB_IN_B16_O)
);
MuxWrapper_1_1 WIRE_SB_T4_WEST_SB_IN_B1 (
    .I(SB_T4_WEST_SB_IN_B1),
    .O(WIRE_SB_T4_WEST_SB_IN_B1_O)
);
MuxWrapper_1_16 WIRE_SB_T4_WEST_SB_IN_B16 (
    .I(SB_T4_WEST_SB_IN_B16),
    .O(WIRE_SB_T4_WEST_SB_IN_B16_O)
);
corebit_and and_inst0 (
    .in0(coreir_eq_16_inst0_out),
    .in1(config_read[0]),
    .out(and_inst0_out)
);
corebit_and and_inst1 (
    .in0(coreir_eq_16_inst0_out),
    .in1(config_write[0]),
    .out(and_inst1_out)
);
coreir_const #(
    .value(8'h00),
    .width(8)
) const_0_8 (
    .out(const_0_8_out)
);
coreir_const #(
    .value(9'h1ff),
    .width(9)
) const_511_9 (
    .out(const_511_9_out)
);
coreir_eq #(
    .width(16)
) coreir_eq_16_inst0 (
    .in0(tile_id),
    .in1(self_config_config_addr_out[15:0]),
    .out(coreir_eq_16_inst0_out)
);
coreir_or #(
    .width(32)
) read_config_data_or_inst0 (
    .in0(read_data_mux_O),
    .in1(read_config_data_in),
    .out(read_config_data_or_inst0_out)
);
MuxWithDefaultWrapper_9_32_8_0 read_data_mux (
    .EN(and_inst0_out),
    .I_0(PE_inst0_read_config_data),
    .I_1(CB_inputs0_read_config_data),
    .I_2(CB_inputs1_read_config_data),
    .I_3(CB_inputs2_read_config_data),
    .I_4(CB_inputs3_read_config_data),
    .I_5(CB_inputs4_read_config_data),
    .I_6(CB_inputs5_read_config_data),
    .I_7(SB_ID0_5TRACKS_B1_PE_read_config_data),
    .I_8(SB_ID0_5TRACKS_B16_PE_read_config_data),
    .O(read_data_mux_O),
    .S(read_data_mux_S_in)
);
mantle_wire__typeBitIn8 read_data_mux_S (
    .in(read_data_mux_S_in),
    .out(self_config_config_addr_out[23:16])
);
mantle_wire__typeBit32 self_config_config_addr (
    .in(config_config_addr),
    .out(self_config_config_addr_out)
);
assign SB_T0_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T0_EAST_SB_OUT_B1;
assign SB_T0_EAST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T0_EAST_SB_OUT_B16;
assign SB_T0_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T0_NORTH_SB_OUT_B1;
assign SB_T0_NORTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T0_NORTH_SB_OUT_B16;
assign SB_T0_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T0_SOUTH_SB_OUT_B1;
assign SB_T0_SOUTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T0_SOUTH_SB_OUT_B16;
assign SB_T0_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T0_WEST_SB_OUT_B1;
assign SB_T0_WEST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T0_WEST_SB_OUT_B16;
assign SB_T1_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T1_EAST_SB_OUT_B1;
assign SB_T1_EAST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T1_EAST_SB_OUT_B16;
assign SB_T1_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T1_NORTH_SB_OUT_B1;
assign SB_T1_NORTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T1_NORTH_SB_OUT_B16;
assign SB_T1_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T1_SOUTH_SB_OUT_B1;
assign SB_T1_SOUTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T1_SOUTH_SB_OUT_B16;
assign SB_T1_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T1_WEST_SB_OUT_B1;
assign SB_T1_WEST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T1_WEST_SB_OUT_B16;
assign SB_T2_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T2_EAST_SB_OUT_B1;
assign SB_T2_EAST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T2_EAST_SB_OUT_B16;
assign SB_T2_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T2_NORTH_SB_OUT_B1;
assign SB_T2_NORTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T2_NORTH_SB_OUT_B16;
assign SB_T2_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T2_SOUTH_SB_OUT_B1;
assign SB_T2_SOUTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T2_SOUTH_SB_OUT_B16;
assign SB_T2_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T2_WEST_SB_OUT_B1;
assign SB_T2_WEST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T2_WEST_SB_OUT_B16;
assign SB_T3_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T3_EAST_SB_OUT_B1;
assign SB_T3_EAST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T3_EAST_SB_OUT_B16;
assign SB_T3_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T3_NORTH_SB_OUT_B1;
assign SB_T3_NORTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T3_NORTH_SB_OUT_B16;
assign SB_T3_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T3_SOUTH_SB_OUT_B1;
assign SB_T3_SOUTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T3_SOUTH_SB_OUT_B16;
assign SB_T3_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T3_WEST_SB_OUT_B1;
assign SB_T3_WEST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T3_WEST_SB_OUT_B16;
assign SB_T4_EAST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T4_EAST_SB_OUT_B1;
assign SB_T4_EAST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T4_EAST_SB_OUT_B16;
assign SB_T4_NORTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T4_NORTH_SB_OUT_B1;
assign SB_T4_NORTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T4_NORTH_SB_OUT_B16;
assign SB_T4_SOUTH_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T4_SOUTH_SB_OUT_B1;
assign SB_T4_SOUTH_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T4_SOUTH_SB_OUT_B16;
assign SB_T4_WEST_SB_OUT_B1 = SB_ID0_5TRACKS_B1_PE_SB_T4_WEST_SB_OUT_B1;
assign SB_T4_WEST_SB_OUT_B16 = SB_ID0_5TRACKS_B16_PE_SB_T4_WEST_SB_OUT_B16;
assign clk_out = clk_pass_through;
assign clk_pass_through_out_bot = clk_pass_through;
assign clk_pass_through_out_right = clk_pass_through;
assign config_out_config_addr = config_config_addr;
assign config_out_config_data = config_config_data;
assign config_out_read = config_read;
assign config_out_write = config_write;
assign hi = const_511_9_out;
assign lo = const_0_8_out;
assign read_config_data = read_config_data_or_inst0_out;
assign reset_out = reset;
assign stall_out = stall;
endmodule

module Interconnect (
    input clk,
    input [31:0] config_0_config_addr,
    input [31:0] config_0_config_data,
    input [0:0] config_0_read,
    input [0:0] config_0_write,
    input [31:0] config_10_config_addr,
    input [31:0] config_10_config_data,
    input [0:0] config_10_read,
    input [0:0] config_10_write,
    input [31:0] config_11_config_addr,
    input [31:0] config_11_config_data,
    input [0:0] config_11_read,
    input [0:0] config_11_write,
    input [31:0] config_12_config_addr,
    input [31:0] config_12_config_data,
    input [0:0] config_12_read,
    input [0:0] config_12_write,
    input [31:0] config_13_config_addr,
    input [31:0] config_13_config_data,
    input [0:0] config_13_read,
    input [0:0] config_13_write,
    input [31:0] config_14_config_addr,
    input [31:0] config_14_config_data,
    input [0:0] config_14_read,
    input [0:0] config_14_write,
    input [31:0] config_15_config_addr,
    input [31:0] config_15_config_data,
    input [0:0] config_15_read,
    input [0:0] config_15_write,
    input [31:0] config_1_config_addr,
    input [31:0] config_1_config_data,
    input [0:0] config_1_read,
    input [0:0] config_1_write,
    input [31:0] config_2_config_addr,
    input [31:0] config_2_config_data,
    input [0:0] config_2_read,
    input [0:0] config_2_write,
    input [31:0] config_3_config_addr,
    input [31:0] config_3_config_data,
    input [0:0] config_3_read,
    input [0:0] config_3_write,
    input [31:0] config_4_config_addr,
    input [31:0] config_4_config_data,
    input [0:0] config_4_read,
    input [0:0] config_4_write,
    input [31:0] config_5_config_addr,
    input [31:0] config_5_config_data,
    input [0:0] config_5_read,
    input [0:0] config_5_write,
    input [31:0] config_6_config_addr,
    input [31:0] config_6_config_data,
    input [0:0] config_6_read,
    input [0:0] config_6_write,
    input [31:0] config_7_config_addr,
    input [31:0] config_7_config_data,
    input [0:0] config_7_read,
    input [0:0] config_7_write,
    input [31:0] config_8_config_addr,
    input [31:0] config_8_config_data,
    input [0:0] config_8_read,
    input [0:0] config_8_write,
    input [31:0] config_9_config_addr,
    input [31:0] config_9_config_data,
    input [0:0] config_9_read,
    input [0:0] config_9_write,
    input [15:0] glb2io_16_X00_Y00,
    input [15:0] glb2io_16_X01_Y00,
    input [15:0] glb2io_16_X02_Y00,
    input [15:0] glb2io_16_X03_Y00,
    input [15:0] glb2io_16_X04_Y00,
    input [15:0] glb2io_16_X05_Y00,
    input [15:0] glb2io_16_X06_Y00,
    input [15:0] glb2io_16_X07_Y00,
    input [15:0] glb2io_16_X08_Y00,
    input [15:0] glb2io_16_X09_Y00,
    input [15:0] glb2io_16_X0A_Y00,
    input [15:0] glb2io_16_X0B_Y00,
    input [15:0] glb2io_16_X0C_Y00,
    input [15:0] glb2io_16_X0D_Y00,
    input [15:0] glb2io_16_X0E_Y00,
    input [15:0] glb2io_16_X0F_Y00,
    input [0:0] glb2io_1_X00_Y00,
    input [0:0] glb2io_1_X01_Y00,
    input [0:0] glb2io_1_X02_Y00,
    input [0:0] glb2io_1_X03_Y00,
    input [0:0] glb2io_1_X04_Y00,
    input [0:0] glb2io_1_X05_Y00,
    input [0:0] glb2io_1_X06_Y00,
    input [0:0] glb2io_1_X07_Y00,
    input [0:0] glb2io_1_X08_Y00,
    input [0:0] glb2io_1_X09_Y00,
    input [0:0] glb2io_1_X0A_Y00,
    input [0:0] glb2io_1_X0B_Y00,
    input [0:0] glb2io_1_X0C_Y00,
    input [0:0] glb2io_1_X0D_Y00,
    input [0:0] glb2io_1_X0E_Y00,
    input [0:0] glb2io_1_X0F_Y00,
    output [15:0] io2glb_16_X00_Y00,
    output [15:0] io2glb_16_X01_Y00,
    output [15:0] io2glb_16_X02_Y00,
    output [15:0] io2glb_16_X03_Y00,
    output [15:0] io2glb_16_X04_Y00,
    output [15:0] io2glb_16_X05_Y00,
    output [15:0] io2glb_16_X06_Y00,
    output [15:0] io2glb_16_X07_Y00,
    output [15:0] io2glb_16_X08_Y00,
    output [15:0] io2glb_16_X09_Y00,
    output [15:0] io2glb_16_X0A_Y00,
    output [15:0] io2glb_16_X0B_Y00,
    output [15:0] io2glb_16_X0C_Y00,
    output [15:0] io2glb_16_X0D_Y00,
    output [15:0] io2glb_16_X0E_Y00,
    output [15:0] io2glb_16_X0F_Y00,
    output [0:0] io2glb_1_X00_Y00,
    output [0:0] io2glb_1_X01_Y00,
    output [0:0] io2glb_1_X02_Y00,
    output [0:0] io2glb_1_X03_Y00,
    output [0:0] io2glb_1_X04_Y00,
    output [0:0] io2glb_1_X05_Y00,
    output [0:0] io2glb_1_X06_Y00,
    output [0:0] io2glb_1_X07_Y00,
    output [0:0] io2glb_1_X08_Y00,
    output [0:0] io2glb_1_X09_Y00,
    output [0:0] io2glb_1_X0A_Y00,
    output [0:0] io2glb_1_X0B_Y00,
    output [0:0] io2glb_1_X0C_Y00,
    output [0:0] io2glb_1_X0D_Y00,
    output [0:0] io2glb_1_X0E_Y00,
    output [0:0] io2glb_1_X0F_Y00,
    output [31:0] read_config_data,
    input reset,
    input [15:0] stall
);
wire [31:0] ConfigPipeStage_inst0_config_out_config_addr;
wire [31:0] ConfigPipeStage_inst0_config_out_config_data;
wire [0:0] ConfigPipeStage_inst0_config_out_read;
wire [0:0] ConfigPipeStage_inst0_config_out_write;
wire [31:0] ConfigPipeStage_inst1_config_out_config_addr;
wire [31:0] ConfigPipeStage_inst1_config_out_config_data;
wire [0:0] ConfigPipeStage_inst1_config_out_read;
wire [0:0] ConfigPipeStage_inst1_config_out_write;
wire [31:0] ConfigPipeStage_inst10_config_out_config_addr;
wire [31:0] ConfigPipeStage_inst10_config_out_config_data;
wire [0:0] ConfigPipeStage_inst10_config_out_read;
wire [0:0] ConfigPipeStage_inst10_config_out_write;
wire [31:0] ConfigPipeStage_inst11_config_out_config_addr;
wire [31:0] ConfigPipeStage_inst11_config_out_config_data;
wire [0:0] ConfigPipeStage_inst11_config_out_read;
wire [0:0] ConfigPipeStage_inst11_config_out_write;
wire [31:0] ConfigPipeStage_inst12_config_out_config_addr;
wire [31:0] ConfigPipeStage_inst12_config_out_config_data;
wire [0:0] ConfigPipeStage_inst12_config_out_read;
wire [0:0] ConfigPipeStage_inst12_config_out_write;
wire [31:0] ConfigPipeStage_inst13_config_out_config_addr;
wire [31:0] ConfigPipeStage_inst13_config_out_config_data;
wire [0:0] ConfigPipeStage_inst13_config_out_read;
wire [0:0] ConfigPipeStage_inst13_config_out_write;
wire [31:0] ConfigPipeStage_inst14_config_out_config_addr;
wire [31:0] ConfigPipeStage_inst14_config_out_config_data;
wire [0:0] ConfigPipeStage_inst14_config_out_read;
wire [0:0] ConfigPipeStage_inst14_config_out_write;
wire [31:0] ConfigPipeStage_inst15_config_out_config_addr;
wire [31:0] ConfigPipeStage_inst15_config_out_config_data;
wire [0:0] ConfigPipeStage_inst15_config_out_read;
wire [0:0] ConfigPipeStage_inst15_config_out_write;
wire [31:0] ConfigPipeStage_inst2_config_out_config_addr;
wire [31:0] ConfigPipeStage_inst2_config_out_config_data;
wire [0:0] ConfigPipeStage_inst2_config_out_read;
wire [0:0] ConfigPipeStage_inst2_config_out_write;
wire [31:0] ConfigPipeStage_inst3_config_out_config_addr;
wire [31:0] ConfigPipeStage_inst3_config_out_config_data;
wire [0:0] ConfigPipeStage_inst3_config_out_read;
wire [0:0] ConfigPipeStage_inst3_config_out_write;
wire [31:0] ConfigPipeStage_inst4_config_out_config_addr;
wire [31:0] ConfigPipeStage_inst4_config_out_config_data;
wire [0:0] ConfigPipeStage_inst4_config_out_read;
wire [0:0] ConfigPipeStage_inst4_config_out_write;
wire [31:0] ConfigPipeStage_inst5_config_out_config_addr;
wire [31:0] ConfigPipeStage_inst5_config_out_config_data;
wire [0:0] ConfigPipeStage_inst5_config_out_read;
wire [0:0] ConfigPipeStage_inst5_config_out_write;
wire [31:0] ConfigPipeStage_inst6_config_out_config_addr;
wire [31:0] ConfigPipeStage_inst6_config_out_config_data;
wire [0:0] ConfigPipeStage_inst6_config_out_read;
wire [0:0] ConfigPipeStage_inst6_config_out_write;
wire [31:0] ConfigPipeStage_inst7_config_out_config_addr;
wire [31:0] ConfigPipeStage_inst7_config_out_config_data;
wire [0:0] ConfigPipeStage_inst7_config_out_read;
wire [0:0] ConfigPipeStage_inst7_config_out_write;
wire [31:0] ConfigPipeStage_inst8_config_out_config_addr;
wire [31:0] ConfigPipeStage_inst8_config_out_config_data;
wire [0:0] ConfigPipeStage_inst8_config_out_read;
wire [0:0] ConfigPipeStage_inst8_config_out_write;
wire [31:0] ConfigPipeStage_inst9_config_out_config_addr;
wire [31:0] ConfigPipeStage_inst9_config_out_config_data;
wire [0:0] ConfigPipeStage_inst9_config_out_read;
wire [0:0] ConfigPipeStage_inst9_config_out_write;
wire [0:0] Tile_X00_Y00_io2glb_1;
wire [0:0] Tile_X00_Y00_io2f_1;
wire [15:0] Tile_X00_Y00_io2glb_16;
wire [15:0] Tile_X00_Y00_io2f_16;
wire [8:0] Tile_X00_Y00_hi;
wire [7:0] Tile_X00_Y00_lo;
wire [0:0] Tile_X00_Y01_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y01_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y01_SB_T4_WEST_SB_OUT_B16;
wire Tile_X00_Y01_clk_out;
wire Tile_X00_Y01_clk_pass_through_out_bot;
wire Tile_X00_Y01_clk_pass_through_out_right;
wire [31:0] Tile_X00_Y01_config_out_config_addr;
wire [31:0] Tile_X00_Y01_config_out_config_data;
wire [0:0] Tile_X00_Y01_config_out_read;
wire [0:0] Tile_X00_Y01_config_out_write;
wire [8:0] Tile_X00_Y01_hi;
wire [7:0] Tile_X00_Y01_lo_unq1;
wire [31:0] Tile_X00_Y01_read_config_data;
wire Tile_X00_Y01_reset_out;
wire [0:0] Tile_X00_Y01_stall_out;
wire [7:0] Tile_X00_Y01_lo_out;
wire [15:0] Tile_X00_Y01_tile_id_in;
wire [0:0] Tile_X00_Y02_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y02_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y02_SB_T4_WEST_SB_OUT_B16;
wire Tile_X00_Y02_clk_out;
wire Tile_X00_Y02_clk_pass_through_out_bot;
wire Tile_X00_Y02_clk_pass_through_out_right;
wire [31:0] Tile_X00_Y02_config_out_config_addr;
wire [31:0] Tile_X00_Y02_config_out_config_data;
wire [0:0] Tile_X00_Y02_config_out_read;
wire [0:0] Tile_X00_Y02_config_out_write;
wire [8:0] Tile_X00_Y02_hi;
wire [7:0] Tile_X00_Y02_lo_unq1;
wire [31:0] Tile_X00_Y02_read_config_data;
wire Tile_X00_Y02_reset_out;
wire [0:0] Tile_X00_Y02_stall_out;
wire [7:0] Tile_X00_Y02_lo_out;
wire [15:0] Tile_X00_Y02_tile_id_in;
wire [0:0] Tile_X00_Y03_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y03_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y03_SB_T4_WEST_SB_OUT_B16;
wire Tile_X00_Y03_clk_out;
wire Tile_X00_Y03_clk_pass_through_out_bot;
wire Tile_X00_Y03_clk_pass_through_out_right;
wire [31:0] Tile_X00_Y03_config_out_config_addr;
wire [31:0] Tile_X00_Y03_config_out_config_data;
wire [0:0] Tile_X00_Y03_config_out_read;
wire [0:0] Tile_X00_Y03_config_out_write;
wire [8:0] Tile_X00_Y03_hi_unq1;
wire [7:0] Tile_X00_Y03_lo_unq1;
wire [31:0] Tile_X00_Y03_read_config_data;
wire Tile_X00_Y03_reset_out;
wire [0:0] Tile_X00_Y03_stall_out;
wire [8:0] Tile_X00_Y03_hi_out;
wire [7:0] Tile_X00_Y03_lo_out;
wire [15:0] Tile_X00_Y03_tile_id_in;
wire [0:0] Tile_X00_Y04_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y04_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y04_SB_T4_WEST_SB_OUT_B16;
wire Tile_X00_Y04_clk_out;
wire Tile_X00_Y04_clk_pass_through_out_bot;
wire Tile_X00_Y04_clk_pass_through_out_right;
wire [31:0] Tile_X00_Y04_config_out_config_addr;
wire [31:0] Tile_X00_Y04_config_out_config_data;
wire [0:0] Tile_X00_Y04_config_out_read;
wire [0:0] Tile_X00_Y04_config_out_write;
wire [8:0] Tile_X00_Y04_hi;
wire [7:0] Tile_X00_Y04_lo_unq1;
wire [31:0] Tile_X00_Y04_read_config_data;
wire Tile_X00_Y04_reset_out;
wire [0:0] Tile_X00_Y04_stall_out;
wire [7:0] Tile_X00_Y04_lo_out;
wire [15:0] Tile_X00_Y04_tile_id_in;
wire [0:0] Tile_X00_Y05_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y05_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y05_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y05_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y05_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y05_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y05_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y05_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y05_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y05_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y05_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y05_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y05_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y05_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y05_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y05_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y05_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y05_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y05_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y05_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y05_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y05_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y05_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y05_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y05_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y05_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y05_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y05_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y05_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y05_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y05_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y05_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y05_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y05_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y05_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y05_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y05_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y05_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y05_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y05_SB_T4_WEST_SB_OUT_B16;
wire Tile_X00_Y05_clk_out;
wire Tile_X00_Y05_clk_pass_through_out_bot;
wire Tile_X00_Y05_clk_pass_through_out_right;
wire [31:0] Tile_X00_Y05_config_out_config_addr;
wire [31:0] Tile_X00_Y05_config_out_config_data;
wire [0:0] Tile_X00_Y05_config_out_read;
wire [0:0] Tile_X00_Y05_config_out_write;
wire [8:0] Tile_X00_Y05_hi;
wire [7:0] Tile_X00_Y05_lo_unq1;
wire [31:0] Tile_X00_Y05_read_config_data;
wire Tile_X00_Y05_reset_out;
wire [0:0] Tile_X00_Y05_stall_out;
wire [7:0] Tile_X00_Y05_lo_out;
wire [15:0] Tile_X00_Y05_tile_id_in;
wire [0:0] Tile_X00_Y06_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y06_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y06_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y06_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y06_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y06_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y06_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y06_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y06_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y06_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y06_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y06_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y06_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y06_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y06_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y06_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y06_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y06_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y06_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y06_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y06_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y06_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y06_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y06_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y06_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y06_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y06_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y06_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y06_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y06_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y06_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y06_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y06_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y06_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y06_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y06_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y06_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y06_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y06_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y06_SB_T4_WEST_SB_OUT_B16;
wire Tile_X00_Y06_clk_out;
wire Tile_X00_Y06_clk_pass_through_out_bot;
wire Tile_X00_Y06_clk_pass_through_out_right;
wire [31:0] Tile_X00_Y06_config_out_config_addr;
wire [31:0] Tile_X00_Y06_config_out_config_data;
wire [0:0] Tile_X00_Y06_config_out_read;
wire [0:0] Tile_X00_Y06_config_out_write;
wire [8:0] Tile_X00_Y06_hi;
wire [7:0] Tile_X00_Y06_lo_unq1;
wire [31:0] Tile_X00_Y06_read_config_data;
wire Tile_X00_Y06_reset_out;
wire [0:0] Tile_X00_Y06_stall_out;
wire [7:0] Tile_X00_Y06_lo_out;
wire [15:0] Tile_X00_Y06_tile_id_in;
wire [0:0] Tile_X00_Y07_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y07_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y07_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y07_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y07_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y07_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y07_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y07_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y07_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y07_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y07_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y07_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y07_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y07_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y07_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y07_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y07_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y07_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y07_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y07_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y07_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y07_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y07_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y07_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y07_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y07_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y07_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y07_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y07_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y07_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y07_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y07_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y07_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y07_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y07_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y07_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y07_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y07_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y07_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y07_SB_T4_WEST_SB_OUT_B16;
wire Tile_X00_Y07_clk_out;
wire Tile_X00_Y07_clk_pass_through_out_bot;
wire Tile_X00_Y07_clk_pass_through_out_right;
wire [31:0] Tile_X00_Y07_config_out_config_addr;
wire [31:0] Tile_X00_Y07_config_out_config_data;
wire [0:0] Tile_X00_Y07_config_out_read;
wire [0:0] Tile_X00_Y07_config_out_write;
wire [8:0] Tile_X00_Y07_hi_unq1;
wire [7:0] Tile_X00_Y07_lo_unq1;
wire [31:0] Tile_X00_Y07_read_config_data;
wire Tile_X00_Y07_reset_out;
wire [0:0] Tile_X00_Y07_stall_out;
wire [8:0] Tile_X00_Y07_hi_out;
wire [7:0] Tile_X00_Y07_lo_out;
wire [15:0] Tile_X00_Y07_tile_id_in;
wire [0:0] Tile_X00_Y08_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y08_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y08_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y08_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y08_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y08_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y08_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y08_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y08_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y08_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y08_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y08_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y08_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y08_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y08_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y08_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y08_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y08_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y08_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y08_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y08_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y08_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y08_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y08_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y08_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y08_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y08_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y08_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y08_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y08_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y08_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y08_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y08_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y08_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y08_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y08_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y08_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y08_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y08_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y08_SB_T4_WEST_SB_OUT_B16;
wire Tile_X00_Y08_clk_out;
wire Tile_X00_Y08_clk_pass_through_out_bot;
wire Tile_X00_Y08_clk_pass_through_out_right;
wire [31:0] Tile_X00_Y08_config_out_config_addr;
wire [31:0] Tile_X00_Y08_config_out_config_data;
wire [0:0] Tile_X00_Y08_config_out_read;
wire [0:0] Tile_X00_Y08_config_out_write;
wire [8:0] Tile_X00_Y08_hi;
wire [7:0] Tile_X00_Y08_lo_unq1;
wire [31:0] Tile_X00_Y08_read_config_data;
wire Tile_X00_Y08_reset_out;
wire [0:0] Tile_X00_Y08_stall_out;
wire [7:0] Tile_X00_Y08_lo_out;
wire [15:0] Tile_X00_Y08_tile_id_in;
wire [0:0] Tile_X00_Y09_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y09_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y09_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y09_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y09_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y09_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y09_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y09_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y09_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y09_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y09_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y09_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y09_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y09_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y09_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y09_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y09_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y09_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y09_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y09_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y09_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y09_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y09_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y09_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y09_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y09_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y09_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y09_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y09_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y09_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y09_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y09_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y09_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y09_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y09_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y09_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y09_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y09_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y09_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y09_SB_T4_WEST_SB_OUT_B16;
wire Tile_X00_Y09_clk_out;
wire Tile_X00_Y09_clk_pass_through_out_bot;
wire Tile_X00_Y09_clk_pass_through_out_right;
wire [31:0] Tile_X00_Y09_config_out_config_addr;
wire [31:0] Tile_X00_Y09_config_out_config_data;
wire [0:0] Tile_X00_Y09_config_out_read;
wire [0:0] Tile_X00_Y09_config_out_write;
wire [8:0] Tile_X00_Y09_hi;
wire [7:0] Tile_X00_Y09_lo_unq1;
wire [31:0] Tile_X00_Y09_read_config_data;
wire Tile_X00_Y09_reset_out;
wire [0:0] Tile_X00_Y09_stall_out;
wire [7:0] Tile_X00_Y09_lo_out;
wire [15:0] Tile_X00_Y09_tile_id_in;
wire [0:0] Tile_X00_Y0A_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0A_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0A_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0A_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0A_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0A_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0A_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0A_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0A_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0A_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0A_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0A_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0A_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0A_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0A_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0A_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0A_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0A_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0A_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0A_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0A_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0A_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0A_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0A_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0A_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0A_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0A_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0A_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0A_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0A_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0A_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0A_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0A_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0A_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0A_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0A_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0A_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0A_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0A_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0A_SB_T4_WEST_SB_OUT_B16;
wire Tile_X00_Y0A_clk_out;
wire Tile_X00_Y0A_clk_pass_through_out_bot;
wire Tile_X00_Y0A_clk_pass_through_out_right;
wire [31:0] Tile_X00_Y0A_config_out_config_addr;
wire [31:0] Tile_X00_Y0A_config_out_config_data;
wire [0:0] Tile_X00_Y0A_config_out_read;
wire [0:0] Tile_X00_Y0A_config_out_write;
wire [8:0] Tile_X00_Y0A_hi;
wire [7:0] Tile_X00_Y0A_lo_unq1;
wire [31:0] Tile_X00_Y0A_read_config_data;
wire Tile_X00_Y0A_reset_out;
wire [0:0] Tile_X00_Y0A_stall_out;
wire [7:0] Tile_X00_Y0A_lo_out;
wire [15:0] Tile_X00_Y0A_tile_id_in;
wire [0:0] Tile_X00_Y0B_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0B_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0B_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0B_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0B_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0B_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0B_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0B_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0B_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0B_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0B_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0B_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0B_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0B_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0B_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0B_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0B_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0B_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0B_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0B_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0B_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0B_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0B_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0B_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0B_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0B_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0B_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0B_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0B_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0B_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0B_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0B_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0B_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0B_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0B_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0B_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0B_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0B_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0B_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0B_SB_T4_WEST_SB_OUT_B16;
wire Tile_X00_Y0B_clk_out;
wire Tile_X00_Y0B_clk_pass_through_out_bot;
wire Tile_X00_Y0B_clk_pass_through_out_right;
wire [31:0] Tile_X00_Y0B_config_out_config_addr;
wire [31:0] Tile_X00_Y0B_config_out_config_data;
wire [0:0] Tile_X00_Y0B_config_out_read;
wire [0:0] Tile_X00_Y0B_config_out_write;
wire [8:0] Tile_X00_Y0B_hi_unq1;
wire [7:0] Tile_X00_Y0B_lo_unq1;
wire [31:0] Tile_X00_Y0B_read_config_data;
wire Tile_X00_Y0B_reset_out;
wire [0:0] Tile_X00_Y0B_stall_out;
wire [8:0] Tile_X00_Y0B_hi_out;
wire [7:0] Tile_X00_Y0B_lo_out;
wire [15:0] Tile_X00_Y0B_tile_id_in;
wire [0:0] Tile_X00_Y0C_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0C_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0C_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0C_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0C_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0C_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0C_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0C_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0C_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0C_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0C_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0C_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0C_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0C_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0C_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0C_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0C_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0C_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0C_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0C_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0C_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0C_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0C_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0C_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0C_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0C_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0C_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0C_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0C_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0C_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0C_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0C_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0C_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0C_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0C_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0C_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0C_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0C_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0C_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0C_SB_T4_WEST_SB_OUT_B16;
wire Tile_X00_Y0C_clk_out;
wire Tile_X00_Y0C_clk_pass_through_out_bot;
wire Tile_X00_Y0C_clk_pass_through_out_right;
wire [31:0] Tile_X00_Y0C_config_out_config_addr;
wire [31:0] Tile_X00_Y0C_config_out_config_data;
wire [0:0] Tile_X00_Y0C_config_out_read;
wire [0:0] Tile_X00_Y0C_config_out_write;
wire [8:0] Tile_X00_Y0C_hi_unq1;
wire [7:0] Tile_X00_Y0C_lo_unq1;
wire [31:0] Tile_X00_Y0C_read_config_data;
wire Tile_X00_Y0C_reset_out;
wire [0:0] Tile_X00_Y0C_stall_out;
wire [8:0] Tile_X00_Y0C_hi_out;
wire [7:0] Tile_X00_Y0C_lo_out;
wire [15:0] Tile_X00_Y0C_tile_id_in;
wire [0:0] Tile_X00_Y0D_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0D_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0D_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0D_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0D_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0D_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0D_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0D_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0D_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0D_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0D_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0D_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0D_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0D_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0D_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0D_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0D_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0D_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0D_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0D_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0D_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0D_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0D_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0D_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0D_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0D_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0D_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0D_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0D_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0D_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0D_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0D_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0D_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0D_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0D_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0D_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0D_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0D_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0D_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0D_SB_T4_WEST_SB_OUT_B16;
wire Tile_X00_Y0D_clk_out;
wire Tile_X00_Y0D_clk_pass_through_out_bot;
wire Tile_X00_Y0D_clk_pass_through_out_right;
wire [31:0] Tile_X00_Y0D_config_out_config_addr;
wire [31:0] Tile_X00_Y0D_config_out_config_data;
wire [0:0] Tile_X00_Y0D_config_out_read;
wire [0:0] Tile_X00_Y0D_config_out_write;
wire [8:0] Tile_X00_Y0D_hi_unq1;
wire [7:0] Tile_X00_Y0D_lo_unq1;
wire [31:0] Tile_X00_Y0D_read_config_data;
wire Tile_X00_Y0D_reset_out;
wire [0:0] Tile_X00_Y0D_stall_out;
wire [8:0] Tile_X00_Y0D_hi_out;
wire [7:0] Tile_X00_Y0D_lo_out;
wire [15:0] Tile_X00_Y0D_tile_id_in;
wire [0:0] Tile_X00_Y0E_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0E_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0E_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0E_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0E_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0E_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0E_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0E_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0E_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0E_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0E_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0E_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0E_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0E_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0E_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0E_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0E_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0E_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0E_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0E_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0E_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0E_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0E_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0E_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0E_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0E_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0E_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0E_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0E_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0E_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0E_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0E_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0E_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0E_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0E_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0E_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0E_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0E_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0E_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0E_SB_T4_WEST_SB_OUT_B16;
wire Tile_X00_Y0E_clk_out;
wire Tile_X00_Y0E_clk_pass_through_out_bot;
wire Tile_X00_Y0E_clk_pass_through_out_right;
wire [31:0] Tile_X00_Y0E_config_out_config_addr;
wire [31:0] Tile_X00_Y0E_config_out_config_data;
wire [0:0] Tile_X00_Y0E_config_out_read;
wire [0:0] Tile_X00_Y0E_config_out_write;
wire [8:0] Tile_X00_Y0E_hi_unq1;
wire [7:0] Tile_X00_Y0E_lo_unq1;
wire [31:0] Tile_X00_Y0E_read_config_data;
wire Tile_X00_Y0E_reset_out;
wire [0:0] Tile_X00_Y0E_stall_out;
wire [8:0] Tile_X00_Y0E_hi_out;
wire [7:0] Tile_X00_Y0E_lo_out;
wire [15:0] Tile_X00_Y0E_tile_id_in;
wire [0:0] Tile_X00_Y0F_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0F_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0F_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0F_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0F_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0F_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0F_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0F_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0F_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0F_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0F_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0F_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0F_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0F_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0F_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0F_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0F_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0F_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0F_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0F_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0F_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0F_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0F_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0F_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0F_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0F_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0F_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0F_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0F_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0F_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0F_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0F_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0F_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0F_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y0F_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0F_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0F_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y0F_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y0F_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y0F_SB_T4_WEST_SB_OUT_B16;
wire Tile_X00_Y0F_clk_out;
wire Tile_X00_Y0F_clk_pass_through_out_bot;
wire Tile_X00_Y0F_clk_pass_through_out_right;
wire [31:0] Tile_X00_Y0F_config_out_config_addr;
wire [31:0] Tile_X00_Y0F_config_out_config_data;
wire [0:0] Tile_X00_Y0F_config_out_read;
wire [0:0] Tile_X00_Y0F_config_out_write;
wire [8:0] Tile_X00_Y0F_hi_unq1;
wire [7:0] Tile_X00_Y0F_lo_unq1;
wire [31:0] Tile_X00_Y0F_read_config_data;
wire Tile_X00_Y0F_reset_out;
wire [0:0] Tile_X00_Y0F_stall_out;
wire [8:0] Tile_X00_Y0F_hi_out;
wire [7:0] Tile_X00_Y0F_lo_out;
wire [15:0] Tile_X00_Y0F_tile_id_in;
wire [0:0] Tile_X00_Y10_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y10_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y10_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y10_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y10_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y10_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y10_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y10_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y10_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y10_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y10_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y10_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y10_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y10_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y10_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y10_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y10_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y10_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y10_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y10_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y10_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y10_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y10_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y10_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y10_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y10_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y10_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y10_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y10_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y10_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y10_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y10_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X00_Y10_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X00_Y10_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X00_Y10_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y10_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y10_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X00_Y10_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X00_Y10_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X00_Y10_SB_T4_WEST_SB_OUT_B16;
wire Tile_X00_Y10_clk_out;
wire Tile_X00_Y10_clk_pass_through_out_bot;
wire Tile_X00_Y10_clk_pass_through_out_right;
wire [31:0] Tile_X00_Y10_config_out_config_addr;
wire [31:0] Tile_X00_Y10_config_out_config_data;
wire [0:0] Tile_X00_Y10_config_out_read;
wire [0:0] Tile_X00_Y10_config_out_write;
wire [8:0] Tile_X00_Y10_hi;
wire [7:0] Tile_X00_Y10_lo_unq1;
wire [31:0] Tile_X00_Y10_read_config_data;
wire Tile_X00_Y10_reset_out;
wire [0:0] Tile_X00_Y10_stall_out;
wire [7:0] Tile_X00_Y10_lo_out;
wire [15:0] Tile_X00_Y10_tile_id_in;
wire [0:0] Tile_X01_Y00_io2glb_1;
wire [0:0] Tile_X01_Y00_io2f_1;
wire [15:0] Tile_X01_Y00_io2glb_16;
wire [15:0] Tile_X01_Y00_io2f_16;
wire [8:0] Tile_X01_Y00_hi;
wire [7:0] Tile_X01_Y00_lo;
wire [0:0] Tile_X01_Y01_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y01_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y01_SB_T4_WEST_SB_OUT_B16;
wire Tile_X01_Y01_clk_out;
wire Tile_X01_Y01_clk_pass_through_out_bot;
wire Tile_X01_Y01_clk_pass_through_out_right;
wire [31:0] Tile_X01_Y01_config_out_config_addr;
wire [31:0] Tile_X01_Y01_config_out_config_data;
wire [0:0] Tile_X01_Y01_config_out_read;
wire [0:0] Tile_X01_Y01_config_out_write;
wire [8:0] Tile_X01_Y01_hi;
wire [7:0] Tile_X01_Y01_lo_unq1;
wire [31:0] Tile_X01_Y01_read_config_data;
wire Tile_X01_Y01_reset_out;
wire [0:0] Tile_X01_Y01_stall_out;
wire [7:0] Tile_X01_Y01_lo_out;
wire [15:0] Tile_X01_Y01_tile_id_in;
wire [0:0] Tile_X01_Y02_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y02_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y02_SB_T4_WEST_SB_OUT_B16;
wire Tile_X01_Y02_clk_out;
wire Tile_X01_Y02_clk_pass_through_out_bot;
wire Tile_X01_Y02_clk_pass_through_out_right;
wire [31:0] Tile_X01_Y02_config_out_config_addr;
wire [31:0] Tile_X01_Y02_config_out_config_data;
wire [0:0] Tile_X01_Y02_config_out_read;
wire [0:0] Tile_X01_Y02_config_out_write;
wire [8:0] Tile_X01_Y02_hi;
wire [7:0] Tile_X01_Y02_lo_unq1;
wire [31:0] Tile_X01_Y02_read_config_data;
wire Tile_X01_Y02_reset_out;
wire [0:0] Tile_X01_Y02_stall_out;
wire [7:0] Tile_X01_Y02_lo_out;
wire [15:0] Tile_X01_Y02_tile_id_in;
wire [0:0] Tile_X01_Y03_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y03_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y03_SB_T4_WEST_SB_OUT_B16;
wire Tile_X01_Y03_clk_out;
wire Tile_X01_Y03_clk_pass_through_out_bot;
wire Tile_X01_Y03_clk_pass_through_out_right;
wire [31:0] Tile_X01_Y03_config_out_config_addr;
wire [31:0] Tile_X01_Y03_config_out_config_data;
wire [0:0] Tile_X01_Y03_config_out_read;
wire [0:0] Tile_X01_Y03_config_out_write;
wire [8:0] Tile_X01_Y03_hi_unq1;
wire [7:0] Tile_X01_Y03_lo_unq1;
wire [31:0] Tile_X01_Y03_read_config_data;
wire Tile_X01_Y03_reset_out;
wire [0:0] Tile_X01_Y03_stall_out;
wire [8:0] Tile_X01_Y03_hi_out;
wire [7:0] Tile_X01_Y03_lo_out;
wire [15:0] Tile_X01_Y03_tile_id_in;
wire [0:0] Tile_X01_Y04_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y04_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y04_SB_T4_WEST_SB_OUT_B16;
wire Tile_X01_Y04_clk_out;
wire Tile_X01_Y04_clk_pass_through_out_bot;
wire Tile_X01_Y04_clk_pass_through_out_right;
wire [31:0] Tile_X01_Y04_config_out_config_addr;
wire [31:0] Tile_X01_Y04_config_out_config_data;
wire [0:0] Tile_X01_Y04_config_out_read;
wire [0:0] Tile_X01_Y04_config_out_write;
wire [8:0] Tile_X01_Y04_hi;
wire [7:0] Tile_X01_Y04_lo_unq1;
wire [31:0] Tile_X01_Y04_read_config_data;
wire Tile_X01_Y04_reset_out;
wire [0:0] Tile_X01_Y04_stall_out;
wire [7:0] Tile_X01_Y04_lo_out;
wire [15:0] Tile_X01_Y04_tile_id_in;
wire [0:0] Tile_X01_Y05_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y05_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y05_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y05_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y05_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y05_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y05_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y05_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y05_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y05_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y05_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y05_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y05_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y05_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y05_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y05_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y05_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y05_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y05_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y05_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y05_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y05_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y05_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y05_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y05_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y05_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y05_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y05_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y05_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y05_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y05_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y05_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y05_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y05_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y05_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y05_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y05_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y05_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y05_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y05_SB_T4_WEST_SB_OUT_B16;
wire Tile_X01_Y05_clk_out;
wire Tile_X01_Y05_clk_pass_through_out_bot;
wire Tile_X01_Y05_clk_pass_through_out_right;
wire [31:0] Tile_X01_Y05_config_out_config_addr;
wire [31:0] Tile_X01_Y05_config_out_config_data;
wire [0:0] Tile_X01_Y05_config_out_read;
wire [0:0] Tile_X01_Y05_config_out_write;
wire [8:0] Tile_X01_Y05_hi;
wire [7:0] Tile_X01_Y05_lo_unq1;
wire [31:0] Tile_X01_Y05_read_config_data;
wire Tile_X01_Y05_reset_out;
wire [0:0] Tile_X01_Y05_stall_out;
wire [7:0] Tile_X01_Y05_lo_out;
wire [15:0] Tile_X01_Y05_tile_id_in;
wire [0:0] Tile_X01_Y06_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y06_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y06_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y06_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y06_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y06_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y06_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y06_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y06_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y06_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y06_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y06_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y06_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y06_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y06_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y06_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y06_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y06_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y06_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y06_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y06_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y06_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y06_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y06_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y06_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y06_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y06_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y06_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y06_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y06_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y06_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y06_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y06_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y06_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y06_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y06_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y06_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y06_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y06_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y06_SB_T4_WEST_SB_OUT_B16;
wire Tile_X01_Y06_clk_out;
wire Tile_X01_Y06_clk_pass_through_out_bot;
wire Tile_X01_Y06_clk_pass_through_out_right;
wire [31:0] Tile_X01_Y06_config_out_config_addr;
wire [31:0] Tile_X01_Y06_config_out_config_data;
wire [0:0] Tile_X01_Y06_config_out_read;
wire [0:0] Tile_X01_Y06_config_out_write;
wire [8:0] Tile_X01_Y06_hi;
wire [7:0] Tile_X01_Y06_lo_unq1;
wire [31:0] Tile_X01_Y06_read_config_data;
wire Tile_X01_Y06_reset_out;
wire [0:0] Tile_X01_Y06_stall_out;
wire [7:0] Tile_X01_Y06_lo_out;
wire [15:0] Tile_X01_Y06_tile_id_in;
wire [0:0] Tile_X01_Y07_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y07_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y07_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y07_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y07_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y07_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y07_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y07_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y07_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y07_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y07_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y07_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y07_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y07_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y07_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y07_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y07_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y07_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y07_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y07_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y07_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y07_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y07_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y07_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y07_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y07_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y07_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y07_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y07_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y07_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y07_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y07_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y07_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y07_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y07_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y07_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y07_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y07_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y07_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y07_SB_T4_WEST_SB_OUT_B16;
wire Tile_X01_Y07_clk_out;
wire Tile_X01_Y07_clk_pass_through_out_bot;
wire Tile_X01_Y07_clk_pass_through_out_right;
wire [31:0] Tile_X01_Y07_config_out_config_addr;
wire [31:0] Tile_X01_Y07_config_out_config_data;
wire [0:0] Tile_X01_Y07_config_out_read;
wire [0:0] Tile_X01_Y07_config_out_write;
wire [8:0] Tile_X01_Y07_hi_unq1;
wire [7:0] Tile_X01_Y07_lo_unq1;
wire [31:0] Tile_X01_Y07_read_config_data;
wire Tile_X01_Y07_reset_out;
wire [0:0] Tile_X01_Y07_stall_out;
wire [8:0] Tile_X01_Y07_hi_out;
wire [7:0] Tile_X01_Y07_lo_out;
wire [15:0] Tile_X01_Y07_tile_id_in;
wire [0:0] Tile_X01_Y08_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y08_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y08_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y08_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y08_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y08_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y08_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y08_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y08_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y08_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y08_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y08_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y08_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y08_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y08_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y08_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y08_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y08_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y08_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y08_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y08_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y08_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y08_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y08_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y08_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y08_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y08_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y08_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y08_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y08_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y08_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y08_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y08_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y08_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y08_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y08_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y08_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y08_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y08_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y08_SB_T4_WEST_SB_OUT_B16;
wire Tile_X01_Y08_clk_out;
wire Tile_X01_Y08_clk_pass_through_out_bot;
wire Tile_X01_Y08_clk_pass_through_out_right;
wire [31:0] Tile_X01_Y08_config_out_config_addr;
wire [31:0] Tile_X01_Y08_config_out_config_data;
wire [0:0] Tile_X01_Y08_config_out_read;
wire [0:0] Tile_X01_Y08_config_out_write;
wire [8:0] Tile_X01_Y08_hi;
wire [7:0] Tile_X01_Y08_lo_unq1;
wire [31:0] Tile_X01_Y08_read_config_data;
wire Tile_X01_Y08_reset_out;
wire [0:0] Tile_X01_Y08_stall_out;
wire [7:0] Tile_X01_Y08_lo_out;
wire [15:0] Tile_X01_Y08_tile_id_in;
wire [0:0] Tile_X01_Y09_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y09_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y09_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y09_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y09_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y09_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y09_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y09_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y09_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y09_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y09_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y09_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y09_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y09_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y09_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y09_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y09_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y09_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y09_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y09_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y09_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y09_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y09_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y09_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y09_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y09_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y09_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y09_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y09_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y09_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y09_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y09_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y09_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y09_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y09_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y09_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y09_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y09_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y09_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y09_SB_T4_WEST_SB_OUT_B16;
wire Tile_X01_Y09_clk_out;
wire Tile_X01_Y09_clk_pass_through_out_bot;
wire Tile_X01_Y09_clk_pass_through_out_right;
wire [31:0] Tile_X01_Y09_config_out_config_addr;
wire [31:0] Tile_X01_Y09_config_out_config_data;
wire [0:0] Tile_X01_Y09_config_out_read;
wire [0:0] Tile_X01_Y09_config_out_write;
wire [8:0] Tile_X01_Y09_hi;
wire [7:0] Tile_X01_Y09_lo_unq1;
wire [31:0] Tile_X01_Y09_read_config_data;
wire Tile_X01_Y09_reset_out;
wire [0:0] Tile_X01_Y09_stall_out;
wire [7:0] Tile_X01_Y09_lo_out;
wire [15:0] Tile_X01_Y09_tile_id_in;
wire [0:0] Tile_X01_Y0A_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0A_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0A_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0A_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0A_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0A_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0A_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0A_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0A_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0A_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0A_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0A_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0A_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0A_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0A_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0A_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0A_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0A_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0A_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0A_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0A_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0A_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0A_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0A_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0A_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0A_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0A_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0A_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0A_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0A_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0A_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0A_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0A_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0A_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0A_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0A_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0A_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0A_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0A_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0A_SB_T4_WEST_SB_OUT_B16;
wire Tile_X01_Y0A_clk_out;
wire Tile_X01_Y0A_clk_pass_through_out_bot;
wire Tile_X01_Y0A_clk_pass_through_out_right;
wire [31:0] Tile_X01_Y0A_config_out_config_addr;
wire [31:0] Tile_X01_Y0A_config_out_config_data;
wire [0:0] Tile_X01_Y0A_config_out_read;
wire [0:0] Tile_X01_Y0A_config_out_write;
wire [8:0] Tile_X01_Y0A_hi;
wire [7:0] Tile_X01_Y0A_lo_unq1;
wire [31:0] Tile_X01_Y0A_read_config_data;
wire Tile_X01_Y0A_reset_out;
wire [0:0] Tile_X01_Y0A_stall_out;
wire [7:0] Tile_X01_Y0A_lo_out;
wire [15:0] Tile_X01_Y0A_tile_id_in;
wire [0:0] Tile_X01_Y0B_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0B_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0B_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0B_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0B_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0B_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0B_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0B_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0B_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0B_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0B_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0B_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0B_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0B_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0B_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0B_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0B_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0B_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0B_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0B_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0B_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0B_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0B_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0B_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0B_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0B_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0B_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0B_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0B_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0B_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0B_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0B_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0B_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0B_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0B_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0B_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0B_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0B_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0B_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0B_SB_T4_WEST_SB_OUT_B16;
wire Tile_X01_Y0B_clk_out;
wire Tile_X01_Y0B_clk_pass_through_out_bot;
wire Tile_X01_Y0B_clk_pass_through_out_right;
wire [31:0] Tile_X01_Y0B_config_out_config_addr;
wire [31:0] Tile_X01_Y0B_config_out_config_data;
wire [0:0] Tile_X01_Y0B_config_out_read;
wire [0:0] Tile_X01_Y0B_config_out_write;
wire [8:0] Tile_X01_Y0B_hi_unq1;
wire [7:0] Tile_X01_Y0B_lo_unq1;
wire [31:0] Tile_X01_Y0B_read_config_data;
wire Tile_X01_Y0B_reset_out;
wire [0:0] Tile_X01_Y0B_stall_out;
wire [8:0] Tile_X01_Y0B_hi_out;
wire [7:0] Tile_X01_Y0B_lo_out;
wire [15:0] Tile_X01_Y0B_tile_id_in;
wire [0:0] Tile_X01_Y0C_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0C_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0C_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0C_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0C_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0C_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0C_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0C_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0C_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0C_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0C_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0C_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0C_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0C_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0C_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0C_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0C_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0C_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0C_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0C_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0C_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0C_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0C_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0C_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0C_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0C_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0C_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0C_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0C_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0C_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0C_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0C_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0C_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0C_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0C_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0C_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0C_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0C_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0C_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0C_SB_T4_WEST_SB_OUT_B16;
wire Tile_X01_Y0C_clk_out;
wire Tile_X01_Y0C_clk_pass_through_out_bot;
wire Tile_X01_Y0C_clk_pass_through_out_right;
wire [31:0] Tile_X01_Y0C_config_out_config_addr;
wire [31:0] Tile_X01_Y0C_config_out_config_data;
wire [0:0] Tile_X01_Y0C_config_out_read;
wire [0:0] Tile_X01_Y0C_config_out_write;
wire [8:0] Tile_X01_Y0C_hi_unq1;
wire [7:0] Tile_X01_Y0C_lo_unq1;
wire [31:0] Tile_X01_Y0C_read_config_data;
wire Tile_X01_Y0C_reset_out;
wire [0:0] Tile_X01_Y0C_stall_out;
wire [8:0] Tile_X01_Y0C_hi_out;
wire [7:0] Tile_X01_Y0C_lo_out;
wire [15:0] Tile_X01_Y0C_tile_id_in;
wire [0:0] Tile_X01_Y0D_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0D_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0D_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0D_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0D_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0D_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0D_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0D_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0D_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0D_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0D_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0D_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0D_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0D_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0D_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0D_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0D_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0D_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0D_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0D_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0D_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0D_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0D_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0D_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0D_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0D_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0D_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0D_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0D_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0D_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0D_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0D_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0D_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0D_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0D_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0D_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0D_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0D_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0D_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0D_SB_T4_WEST_SB_OUT_B16;
wire Tile_X01_Y0D_clk_out;
wire Tile_X01_Y0D_clk_pass_through_out_bot;
wire Tile_X01_Y0D_clk_pass_through_out_right;
wire [31:0] Tile_X01_Y0D_config_out_config_addr;
wire [31:0] Tile_X01_Y0D_config_out_config_data;
wire [0:0] Tile_X01_Y0D_config_out_read;
wire [0:0] Tile_X01_Y0D_config_out_write;
wire [8:0] Tile_X01_Y0D_hi_unq1;
wire [7:0] Tile_X01_Y0D_lo_unq1;
wire [31:0] Tile_X01_Y0D_read_config_data;
wire Tile_X01_Y0D_reset_out;
wire [0:0] Tile_X01_Y0D_stall_out;
wire [8:0] Tile_X01_Y0D_hi_out;
wire [7:0] Tile_X01_Y0D_lo_out;
wire [15:0] Tile_X01_Y0D_tile_id_in;
wire [0:0] Tile_X01_Y0E_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0E_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0E_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0E_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0E_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0E_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0E_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0E_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0E_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0E_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0E_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0E_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0E_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0E_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0E_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0E_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0E_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0E_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0E_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0E_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0E_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0E_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0E_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0E_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0E_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0E_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0E_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0E_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0E_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0E_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0E_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0E_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0E_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0E_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0E_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0E_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0E_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0E_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0E_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0E_SB_T4_WEST_SB_OUT_B16;
wire Tile_X01_Y0E_clk_out;
wire Tile_X01_Y0E_clk_pass_through_out_bot;
wire Tile_X01_Y0E_clk_pass_through_out_right;
wire [31:0] Tile_X01_Y0E_config_out_config_addr;
wire [31:0] Tile_X01_Y0E_config_out_config_data;
wire [0:0] Tile_X01_Y0E_config_out_read;
wire [0:0] Tile_X01_Y0E_config_out_write;
wire [8:0] Tile_X01_Y0E_hi_unq1;
wire [7:0] Tile_X01_Y0E_lo_unq1;
wire [31:0] Tile_X01_Y0E_read_config_data;
wire Tile_X01_Y0E_reset_out;
wire [0:0] Tile_X01_Y0E_stall_out;
wire [8:0] Tile_X01_Y0E_hi_out;
wire [7:0] Tile_X01_Y0E_lo_out;
wire [15:0] Tile_X01_Y0E_tile_id_in;
wire [0:0] Tile_X01_Y0F_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0F_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0F_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0F_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0F_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0F_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0F_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0F_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0F_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0F_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0F_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0F_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0F_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0F_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0F_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0F_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0F_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0F_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0F_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0F_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0F_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0F_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0F_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0F_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0F_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0F_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0F_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0F_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0F_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0F_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0F_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0F_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0F_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0F_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y0F_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0F_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0F_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y0F_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y0F_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y0F_SB_T4_WEST_SB_OUT_B16;
wire Tile_X01_Y0F_clk_out;
wire Tile_X01_Y0F_clk_pass_through_out_bot;
wire Tile_X01_Y0F_clk_pass_through_out_right;
wire [31:0] Tile_X01_Y0F_config_out_config_addr;
wire [31:0] Tile_X01_Y0F_config_out_config_data;
wire [0:0] Tile_X01_Y0F_config_out_read;
wire [0:0] Tile_X01_Y0F_config_out_write;
wire [8:0] Tile_X01_Y0F_hi_unq1;
wire [7:0] Tile_X01_Y0F_lo_unq1;
wire [31:0] Tile_X01_Y0F_read_config_data;
wire Tile_X01_Y0F_reset_out;
wire [0:0] Tile_X01_Y0F_stall_out;
wire [8:0] Tile_X01_Y0F_hi_out;
wire [7:0] Tile_X01_Y0F_lo_out;
wire [15:0] Tile_X01_Y0F_tile_id_in;
wire [0:0] Tile_X01_Y10_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y10_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y10_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y10_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y10_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y10_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y10_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y10_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y10_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y10_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y10_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y10_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y10_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y10_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y10_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y10_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y10_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y10_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y10_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y10_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y10_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y10_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y10_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y10_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y10_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y10_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y10_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y10_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y10_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y10_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y10_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y10_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X01_Y10_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X01_Y10_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X01_Y10_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y10_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y10_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X01_Y10_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X01_Y10_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X01_Y10_SB_T4_WEST_SB_OUT_B16;
wire Tile_X01_Y10_clk_out;
wire Tile_X01_Y10_clk_pass_through_out_bot;
wire Tile_X01_Y10_clk_pass_through_out_right;
wire [31:0] Tile_X01_Y10_config_out_config_addr;
wire [31:0] Tile_X01_Y10_config_out_config_data;
wire [0:0] Tile_X01_Y10_config_out_read;
wire [0:0] Tile_X01_Y10_config_out_write;
wire [8:0] Tile_X01_Y10_hi;
wire [7:0] Tile_X01_Y10_lo_unq1;
wire [31:0] Tile_X01_Y10_read_config_data;
wire Tile_X01_Y10_reset_out;
wire [0:0] Tile_X01_Y10_stall_out;
wire [7:0] Tile_X01_Y10_lo_out;
wire [15:0] Tile_X01_Y10_tile_id_in;
wire [0:0] Tile_X02_Y00_io2glb_1;
wire [0:0] Tile_X02_Y00_io2f_1;
wire [15:0] Tile_X02_Y00_io2glb_16;
wire [15:0] Tile_X02_Y00_io2f_16;
wire [8:0] Tile_X02_Y00_hi;
wire [7:0] Tile_X02_Y00_lo;
wire [0:0] Tile_X02_Y01_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y01_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y01_SB_T4_WEST_SB_OUT_B16;
wire Tile_X02_Y01_clk_out;
wire Tile_X02_Y01_clk_pass_through_out_bot;
wire Tile_X02_Y01_clk_pass_through_out_right;
wire [31:0] Tile_X02_Y01_config_out_config_addr;
wire [31:0] Tile_X02_Y01_config_out_config_data;
wire [0:0] Tile_X02_Y01_config_out_read;
wire [0:0] Tile_X02_Y01_config_out_write;
wire [8:0] Tile_X02_Y01_hi;
wire [7:0] Tile_X02_Y01_lo_unq1;
wire [31:0] Tile_X02_Y01_read_config_data;
wire Tile_X02_Y01_reset_out;
wire [0:0] Tile_X02_Y01_stall_out;
wire [7:0] Tile_X02_Y01_lo_out;
wire [15:0] Tile_X02_Y01_tile_id_in;
wire [0:0] Tile_X02_Y02_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y02_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y02_SB_T4_WEST_SB_OUT_B16;
wire Tile_X02_Y02_clk_out;
wire Tile_X02_Y02_clk_pass_through_out_bot;
wire Tile_X02_Y02_clk_pass_through_out_right;
wire [31:0] Tile_X02_Y02_config_out_config_addr;
wire [31:0] Tile_X02_Y02_config_out_config_data;
wire [0:0] Tile_X02_Y02_config_out_read;
wire [0:0] Tile_X02_Y02_config_out_write;
wire [8:0] Tile_X02_Y02_hi;
wire [7:0] Tile_X02_Y02_lo_unq1;
wire [31:0] Tile_X02_Y02_read_config_data;
wire Tile_X02_Y02_reset_out;
wire [0:0] Tile_X02_Y02_stall_out;
wire [7:0] Tile_X02_Y02_lo_out;
wire [15:0] Tile_X02_Y02_tile_id_in;
wire [0:0] Tile_X02_Y03_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y03_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y03_SB_T4_WEST_SB_OUT_B16;
wire Tile_X02_Y03_clk_out;
wire Tile_X02_Y03_clk_pass_through_out_bot;
wire Tile_X02_Y03_clk_pass_through_out_right;
wire [31:0] Tile_X02_Y03_config_out_config_addr;
wire [31:0] Tile_X02_Y03_config_out_config_data;
wire [0:0] Tile_X02_Y03_config_out_read;
wire [0:0] Tile_X02_Y03_config_out_write;
wire [8:0] Tile_X02_Y03_hi_unq1;
wire [7:0] Tile_X02_Y03_lo_unq1;
wire [31:0] Tile_X02_Y03_read_config_data;
wire Tile_X02_Y03_reset_out;
wire [0:0] Tile_X02_Y03_stall_out;
wire [8:0] Tile_X02_Y03_hi_out;
wire [7:0] Tile_X02_Y03_lo_out;
wire [15:0] Tile_X02_Y03_tile_id_in;
wire [0:0] Tile_X02_Y04_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y04_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y04_SB_T4_WEST_SB_OUT_B16;
wire Tile_X02_Y04_clk_out;
wire Tile_X02_Y04_clk_pass_through_out_bot;
wire Tile_X02_Y04_clk_pass_through_out_right;
wire [31:0] Tile_X02_Y04_config_out_config_addr;
wire [31:0] Tile_X02_Y04_config_out_config_data;
wire [0:0] Tile_X02_Y04_config_out_read;
wire [0:0] Tile_X02_Y04_config_out_write;
wire [8:0] Tile_X02_Y04_hi;
wire [7:0] Tile_X02_Y04_lo_unq1;
wire [31:0] Tile_X02_Y04_read_config_data;
wire Tile_X02_Y04_reset_out;
wire [0:0] Tile_X02_Y04_stall_out;
wire [7:0] Tile_X02_Y04_lo_out;
wire [15:0] Tile_X02_Y04_tile_id_in;
wire [0:0] Tile_X02_Y05_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y05_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y05_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y05_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y05_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y05_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y05_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y05_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y05_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y05_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y05_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y05_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y05_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y05_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y05_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y05_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y05_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y05_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y05_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y05_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y05_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y05_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y05_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y05_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y05_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y05_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y05_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y05_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y05_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y05_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y05_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y05_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y05_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y05_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y05_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y05_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y05_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y05_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y05_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y05_SB_T4_WEST_SB_OUT_B16;
wire Tile_X02_Y05_clk_out;
wire Tile_X02_Y05_clk_pass_through_out_bot;
wire Tile_X02_Y05_clk_pass_through_out_right;
wire [31:0] Tile_X02_Y05_config_out_config_addr;
wire [31:0] Tile_X02_Y05_config_out_config_data;
wire [0:0] Tile_X02_Y05_config_out_read;
wire [0:0] Tile_X02_Y05_config_out_write;
wire [8:0] Tile_X02_Y05_hi;
wire [7:0] Tile_X02_Y05_lo_unq1;
wire [31:0] Tile_X02_Y05_read_config_data;
wire Tile_X02_Y05_reset_out;
wire [0:0] Tile_X02_Y05_stall_out;
wire [7:0] Tile_X02_Y05_lo_out;
wire [15:0] Tile_X02_Y05_tile_id_in;
wire [0:0] Tile_X02_Y06_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y06_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y06_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y06_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y06_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y06_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y06_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y06_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y06_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y06_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y06_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y06_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y06_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y06_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y06_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y06_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y06_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y06_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y06_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y06_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y06_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y06_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y06_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y06_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y06_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y06_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y06_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y06_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y06_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y06_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y06_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y06_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y06_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y06_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y06_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y06_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y06_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y06_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y06_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y06_SB_T4_WEST_SB_OUT_B16;
wire Tile_X02_Y06_clk_out;
wire Tile_X02_Y06_clk_pass_through_out_bot;
wire Tile_X02_Y06_clk_pass_through_out_right;
wire [31:0] Tile_X02_Y06_config_out_config_addr;
wire [31:0] Tile_X02_Y06_config_out_config_data;
wire [0:0] Tile_X02_Y06_config_out_read;
wire [0:0] Tile_X02_Y06_config_out_write;
wire [8:0] Tile_X02_Y06_hi;
wire [7:0] Tile_X02_Y06_lo_unq1;
wire [31:0] Tile_X02_Y06_read_config_data;
wire Tile_X02_Y06_reset_out;
wire [0:0] Tile_X02_Y06_stall_out;
wire [7:0] Tile_X02_Y06_lo_out;
wire [15:0] Tile_X02_Y06_tile_id_in;
wire [0:0] Tile_X02_Y07_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y07_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y07_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y07_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y07_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y07_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y07_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y07_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y07_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y07_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y07_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y07_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y07_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y07_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y07_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y07_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y07_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y07_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y07_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y07_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y07_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y07_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y07_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y07_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y07_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y07_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y07_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y07_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y07_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y07_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y07_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y07_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y07_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y07_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y07_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y07_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y07_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y07_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y07_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y07_SB_T4_WEST_SB_OUT_B16;
wire Tile_X02_Y07_clk_out;
wire Tile_X02_Y07_clk_pass_through_out_bot;
wire Tile_X02_Y07_clk_pass_through_out_right;
wire [31:0] Tile_X02_Y07_config_out_config_addr;
wire [31:0] Tile_X02_Y07_config_out_config_data;
wire [0:0] Tile_X02_Y07_config_out_read;
wire [0:0] Tile_X02_Y07_config_out_write;
wire [8:0] Tile_X02_Y07_hi_unq1;
wire [7:0] Tile_X02_Y07_lo_unq1;
wire [31:0] Tile_X02_Y07_read_config_data;
wire Tile_X02_Y07_reset_out;
wire [0:0] Tile_X02_Y07_stall_out;
wire [8:0] Tile_X02_Y07_hi_out;
wire [7:0] Tile_X02_Y07_lo_out;
wire [15:0] Tile_X02_Y07_tile_id_in;
wire [0:0] Tile_X02_Y08_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y08_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y08_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y08_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y08_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y08_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y08_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y08_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y08_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y08_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y08_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y08_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y08_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y08_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y08_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y08_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y08_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y08_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y08_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y08_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y08_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y08_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y08_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y08_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y08_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y08_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y08_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y08_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y08_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y08_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y08_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y08_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y08_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y08_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y08_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y08_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y08_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y08_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y08_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y08_SB_T4_WEST_SB_OUT_B16;
wire Tile_X02_Y08_clk_out;
wire Tile_X02_Y08_clk_pass_through_out_bot;
wire Tile_X02_Y08_clk_pass_through_out_right;
wire [31:0] Tile_X02_Y08_config_out_config_addr;
wire [31:0] Tile_X02_Y08_config_out_config_data;
wire [0:0] Tile_X02_Y08_config_out_read;
wire [0:0] Tile_X02_Y08_config_out_write;
wire [8:0] Tile_X02_Y08_hi;
wire [7:0] Tile_X02_Y08_lo_unq1;
wire [31:0] Tile_X02_Y08_read_config_data;
wire Tile_X02_Y08_reset_out;
wire [0:0] Tile_X02_Y08_stall_out;
wire [7:0] Tile_X02_Y08_lo_out;
wire [15:0] Tile_X02_Y08_tile_id_in;
wire [0:0] Tile_X02_Y09_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y09_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y09_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y09_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y09_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y09_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y09_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y09_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y09_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y09_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y09_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y09_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y09_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y09_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y09_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y09_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y09_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y09_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y09_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y09_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y09_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y09_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y09_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y09_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y09_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y09_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y09_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y09_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y09_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y09_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y09_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y09_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y09_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y09_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y09_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y09_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y09_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y09_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y09_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y09_SB_T4_WEST_SB_OUT_B16;
wire Tile_X02_Y09_clk_out;
wire Tile_X02_Y09_clk_pass_through_out_bot;
wire Tile_X02_Y09_clk_pass_through_out_right;
wire [31:0] Tile_X02_Y09_config_out_config_addr;
wire [31:0] Tile_X02_Y09_config_out_config_data;
wire [0:0] Tile_X02_Y09_config_out_read;
wire [0:0] Tile_X02_Y09_config_out_write;
wire [8:0] Tile_X02_Y09_hi;
wire [7:0] Tile_X02_Y09_lo_unq1;
wire [31:0] Tile_X02_Y09_read_config_data;
wire Tile_X02_Y09_reset_out;
wire [0:0] Tile_X02_Y09_stall_out;
wire [7:0] Tile_X02_Y09_lo_out;
wire [15:0] Tile_X02_Y09_tile_id_in;
wire [0:0] Tile_X02_Y0A_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0A_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0A_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0A_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0A_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0A_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0A_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0A_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0A_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0A_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0A_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0A_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0A_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0A_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0A_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0A_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0A_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0A_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0A_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0A_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0A_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0A_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0A_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0A_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0A_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0A_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0A_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0A_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0A_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0A_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0A_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0A_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0A_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0A_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0A_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0A_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0A_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0A_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0A_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0A_SB_T4_WEST_SB_OUT_B16;
wire Tile_X02_Y0A_clk_out;
wire Tile_X02_Y0A_clk_pass_through_out_bot;
wire Tile_X02_Y0A_clk_pass_through_out_right;
wire [31:0] Tile_X02_Y0A_config_out_config_addr;
wire [31:0] Tile_X02_Y0A_config_out_config_data;
wire [0:0] Tile_X02_Y0A_config_out_read;
wire [0:0] Tile_X02_Y0A_config_out_write;
wire [8:0] Tile_X02_Y0A_hi;
wire [7:0] Tile_X02_Y0A_lo_unq1;
wire [31:0] Tile_X02_Y0A_read_config_data;
wire Tile_X02_Y0A_reset_out;
wire [0:0] Tile_X02_Y0A_stall_out;
wire [7:0] Tile_X02_Y0A_lo_out;
wire [15:0] Tile_X02_Y0A_tile_id_in;
wire [0:0] Tile_X02_Y0B_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0B_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0B_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0B_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0B_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0B_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0B_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0B_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0B_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0B_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0B_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0B_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0B_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0B_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0B_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0B_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0B_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0B_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0B_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0B_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0B_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0B_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0B_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0B_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0B_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0B_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0B_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0B_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0B_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0B_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0B_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0B_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0B_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0B_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0B_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0B_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0B_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0B_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0B_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0B_SB_T4_WEST_SB_OUT_B16;
wire Tile_X02_Y0B_clk_out;
wire Tile_X02_Y0B_clk_pass_through_out_bot;
wire Tile_X02_Y0B_clk_pass_through_out_right;
wire [31:0] Tile_X02_Y0B_config_out_config_addr;
wire [31:0] Tile_X02_Y0B_config_out_config_data;
wire [0:0] Tile_X02_Y0B_config_out_read;
wire [0:0] Tile_X02_Y0B_config_out_write;
wire [8:0] Tile_X02_Y0B_hi_unq1;
wire [7:0] Tile_X02_Y0B_lo_unq1;
wire [31:0] Tile_X02_Y0B_read_config_data;
wire Tile_X02_Y0B_reset_out;
wire [0:0] Tile_X02_Y0B_stall_out;
wire [8:0] Tile_X02_Y0B_hi_out;
wire [7:0] Tile_X02_Y0B_lo_out;
wire [15:0] Tile_X02_Y0B_tile_id_in;
wire [0:0] Tile_X02_Y0C_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0C_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0C_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0C_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0C_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0C_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0C_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0C_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0C_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0C_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0C_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0C_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0C_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0C_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0C_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0C_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0C_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0C_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0C_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0C_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0C_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0C_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0C_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0C_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0C_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0C_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0C_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0C_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0C_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0C_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0C_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0C_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0C_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0C_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0C_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0C_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0C_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0C_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0C_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0C_SB_T4_WEST_SB_OUT_B16;
wire Tile_X02_Y0C_clk_out;
wire Tile_X02_Y0C_clk_pass_through_out_bot;
wire Tile_X02_Y0C_clk_pass_through_out_right;
wire [31:0] Tile_X02_Y0C_config_out_config_addr;
wire [31:0] Tile_X02_Y0C_config_out_config_data;
wire [0:0] Tile_X02_Y0C_config_out_read;
wire [0:0] Tile_X02_Y0C_config_out_write;
wire [8:0] Tile_X02_Y0C_hi_unq1;
wire [7:0] Tile_X02_Y0C_lo_unq1;
wire [31:0] Tile_X02_Y0C_read_config_data;
wire Tile_X02_Y0C_reset_out;
wire [0:0] Tile_X02_Y0C_stall_out;
wire [8:0] Tile_X02_Y0C_hi_out;
wire [7:0] Tile_X02_Y0C_lo_out;
wire [15:0] Tile_X02_Y0C_tile_id_in;
wire [0:0] Tile_X02_Y0D_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0D_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0D_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0D_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0D_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0D_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0D_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0D_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0D_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0D_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0D_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0D_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0D_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0D_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0D_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0D_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0D_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0D_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0D_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0D_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0D_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0D_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0D_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0D_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0D_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0D_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0D_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0D_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0D_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0D_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0D_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0D_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0D_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0D_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0D_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0D_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0D_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0D_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0D_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0D_SB_T4_WEST_SB_OUT_B16;
wire Tile_X02_Y0D_clk_out;
wire Tile_X02_Y0D_clk_pass_through_out_bot;
wire Tile_X02_Y0D_clk_pass_through_out_right;
wire [31:0] Tile_X02_Y0D_config_out_config_addr;
wire [31:0] Tile_X02_Y0D_config_out_config_data;
wire [0:0] Tile_X02_Y0D_config_out_read;
wire [0:0] Tile_X02_Y0D_config_out_write;
wire [8:0] Tile_X02_Y0D_hi_unq1;
wire [7:0] Tile_X02_Y0D_lo_unq1;
wire [31:0] Tile_X02_Y0D_read_config_data;
wire Tile_X02_Y0D_reset_out;
wire [0:0] Tile_X02_Y0D_stall_out;
wire [8:0] Tile_X02_Y0D_hi_out;
wire [7:0] Tile_X02_Y0D_lo_out;
wire [15:0] Tile_X02_Y0D_tile_id_in;
wire [0:0] Tile_X02_Y0E_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0E_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0E_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0E_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0E_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0E_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0E_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0E_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0E_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0E_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0E_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0E_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0E_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0E_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0E_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0E_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0E_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0E_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0E_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0E_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0E_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0E_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0E_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0E_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0E_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0E_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0E_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0E_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0E_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0E_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0E_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0E_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0E_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0E_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0E_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0E_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0E_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0E_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0E_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0E_SB_T4_WEST_SB_OUT_B16;
wire Tile_X02_Y0E_clk_out;
wire Tile_X02_Y0E_clk_pass_through_out_bot;
wire Tile_X02_Y0E_clk_pass_through_out_right;
wire [31:0] Tile_X02_Y0E_config_out_config_addr;
wire [31:0] Tile_X02_Y0E_config_out_config_data;
wire [0:0] Tile_X02_Y0E_config_out_read;
wire [0:0] Tile_X02_Y0E_config_out_write;
wire [8:0] Tile_X02_Y0E_hi_unq1;
wire [7:0] Tile_X02_Y0E_lo_unq1;
wire [31:0] Tile_X02_Y0E_read_config_data;
wire Tile_X02_Y0E_reset_out;
wire [0:0] Tile_X02_Y0E_stall_out;
wire [8:0] Tile_X02_Y0E_hi_out;
wire [7:0] Tile_X02_Y0E_lo_out;
wire [15:0] Tile_X02_Y0E_tile_id_in;
wire [0:0] Tile_X02_Y0F_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0F_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0F_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0F_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0F_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0F_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0F_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0F_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0F_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0F_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0F_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0F_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0F_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0F_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0F_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0F_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0F_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0F_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0F_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0F_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0F_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0F_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0F_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0F_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0F_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0F_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0F_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0F_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0F_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0F_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0F_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0F_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0F_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0F_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y0F_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0F_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0F_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y0F_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y0F_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y0F_SB_T4_WEST_SB_OUT_B16;
wire Tile_X02_Y0F_clk_out;
wire Tile_X02_Y0F_clk_pass_through_out_bot;
wire Tile_X02_Y0F_clk_pass_through_out_right;
wire [31:0] Tile_X02_Y0F_config_out_config_addr;
wire [31:0] Tile_X02_Y0F_config_out_config_data;
wire [0:0] Tile_X02_Y0F_config_out_read;
wire [0:0] Tile_X02_Y0F_config_out_write;
wire [8:0] Tile_X02_Y0F_hi_unq1;
wire [7:0] Tile_X02_Y0F_lo_unq1;
wire [31:0] Tile_X02_Y0F_read_config_data;
wire Tile_X02_Y0F_reset_out;
wire [0:0] Tile_X02_Y0F_stall_out;
wire [8:0] Tile_X02_Y0F_hi_out;
wire [7:0] Tile_X02_Y0F_lo_out;
wire [15:0] Tile_X02_Y0F_tile_id_in;
wire [0:0] Tile_X02_Y10_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y10_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y10_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y10_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y10_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y10_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y10_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y10_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y10_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y10_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y10_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y10_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y10_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y10_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y10_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y10_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y10_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y10_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y10_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y10_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y10_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y10_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y10_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y10_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y10_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y10_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y10_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y10_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y10_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y10_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y10_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y10_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X02_Y10_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X02_Y10_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X02_Y10_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y10_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y10_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X02_Y10_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X02_Y10_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X02_Y10_SB_T4_WEST_SB_OUT_B16;
wire Tile_X02_Y10_clk_out;
wire Tile_X02_Y10_clk_pass_through_out_bot;
wire Tile_X02_Y10_clk_pass_through_out_right;
wire [31:0] Tile_X02_Y10_config_out_config_addr;
wire [31:0] Tile_X02_Y10_config_out_config_data;
wire [0:0] Tile_X02_Y10_config_out_read;
wire [0:0] Tile_X02_Y10_config_out_write;
wire [8:0] Tile_X02_Y10_hi;
wire [7:0] Tile_X02_Y10_lo_unq1;
wire [31:0] Tile_X02_Y10_read_config_data;
wire Tile_X02_Y10_reset_out;
wire [0:0] Tile_X02_Y10_stall_out;
wire [7:0] Tile_X02_Y10_lo_out;
wire [15:0] Tile_X02_Y10_tile_id_in;
wire [0:0] Tile_X03_Y00_io2glb_1;
wire [0:0] Tile_X03_Y00_io2f_1;
wire [15:0] Tile_X03_Y00_io2glb_16;
wire [15:0] Tile_X03_Y00_io2f_16;
wire [8:0] Tile_X03_Y00_hi;
wire [7:0] Tile_X03_Y00_lo;
wire [0:0] Tile_X03_Y01_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y01_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y01_SB_T4_WEST_SB_OUT_B16;
wire Tile_X03_Y01_clk_out;
wire [31:0] Tile_X03_Y01_config_out_config_addr;
wire [31:0] Tile_X03_Y01_config_out_config_data;
wire [0:0] Tile_X03_Y01_config_out_read;
wire [0:0] Tile_X03_Y01_config_out_write;
wire [8:0] Tile_X03_Y01_hi_unq1;
wire [7:0] Tile_X03_Y01_lo_unq1;
wire [31:0] Tile_X03_Y01_read_config_data;
wire Tile_X03_Y01_reset_out;
wire [0:0] Tile_X03_Y01_stall_out;
wire [8:0] Tile_X03_Y01_hi_out;
wire [7:0] Tile_X03_Y01_lo_out;
wire [15:0] Tile_X03_Y01_tile_id_in;
wire [0:0] Tile_X03_Y02_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y02_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y02_SB_T4_WEST_SB_OUT_B16;
wire Tile_X03_Y02_clk_out;
wire [31:0] Tile_X03_Y02_config_out_config_addr;
wire [31:0] Tile_X03_Y02_config_out_config_data;
wire [0:0] Tile_X03_Y02_config_out_read;
wire [0:0] Tile_X03_Y02_config_out_write;
wire [8:0] Tile_X03_Y02_hi_unq1;
wire [7:0] Tile_X03_Y02_lo_unq1;
wire [31:0] Tile_X03_Y02_read_config_data;
wire Tile_X03_Y02_reset_out;
wire [0:0] Tile_X03_Y02_stall_out;
wire [8:0] Tile_X03_Y02_hi_out;
wire [7:0] Tile_X03_Y02_lo_out;
wire [15:0] Tile_X03_Y02_tile_id_in;
wire [0:0] Tile_X03_Y03_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y03_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y03_SB_T4_WEST_SB_OUT_B16;
wire Tile_X03_Y03_clk_out;
wire [31:0] Tile_X03_Y03_config_out_config_addr;
wire [31:0] Tile_X03_Y03_config_out_config_data;
wire [0:0] Tile_X03_Y03_config_out_read;
wire [0:0] Tile_X03_Y03_config_out_write;
wire [8:0] Tile_X03_Y03_hi_unq1;
wire [7:0] Tile_X03_Y03_lo_unq1;
wire [31:0] Tile_X03_Y03_read_config_data;
wire Tile_X03_Y03_reset_out;
wire [0:0] Tile_X03_Y03_stall_out;
wire [8:0] Tile_X03_Y03_hi_out;
wire [7:0] Tile_X03_Y03_lo_out;
wire [15:0] Tile_X03_Y03_tile_id_in;
wire [0:0] Tile_X03_Y04_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y04_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y04_SB_T4_WEST_SB_OUT_B16;
wire Tile_X03_Y04_clk_out;
wire [31:0] Tile_X03_Y04_config_out_config_addr;
wire [31:0] Tile_X03_Y04_config_out_config_data;
wire [0:0] Tile_X03_Y04_config_out_read;
wire [0:0] Tile_X03_Y04_config_out_write;
wire [8:0] Tile_X03_Y04_hi_unq1;
wire [7:0] Tile_X03_Y04_lo_unq1;
wire [31:0] Tile_X03_Y04_read_config_data;
wire Tile_X03_Y04_reset_out;
wire [0:0] Tile_X03_Y04_stall_out;
wire [8:0] Tile_X03_Y04_hi_out;
wire [7:0] Tile_X03_Y04_lo_out;
wire [15:0] Tile_X03_Y04_tile_id_in;
wire [0:0] Tile_X03_Y05_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y05_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y05_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y05_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y05_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y05_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y05_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y05_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y05_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y05_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y05_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y05_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y05_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y05_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y05_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y05_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y05_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y05_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y05_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y05_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y05_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y05_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y05_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y05_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y05_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y05_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y05_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y05_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y05_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y05_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y05_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y05_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y05_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y05_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y05_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y05_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y05_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y05_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y05_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y05_SB_T4_WEST_SB_OUT_B16;
wire Tile_X03_Y05_clk_out;
wire [31:0] Tile_X03_Y05_config_out_config_addr;
wire [31:0] Tile_X03_Y05_config_out_config_data;
wire [0:0] Tile_X03_Y05_config_out_read;
wire [0:0] Tile_X03_Y05_config_out_write;
wire [8:0] Tile_X03_Y05_hi_unq1;
wire [7:0] Tile_X03_Y05_lo_unq1;
wire [31:0] Tile_X03_Y05_read_config_data;
wire Tile_X03_Y05_reset_out;
wire [0:0] Tile_X03_Y05_stall_out;
wire [8:0] Tile_X03_Y05_hi_out;
wire [7:0] Tile_X03_Y05_lo_out;
wire [15:0] Tile_X03_Y05_tile_id_in;
wire [0:0] Tile_X03_Y06_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y06_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y06_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y06_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y06_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y06_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y06_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y06_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y06_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y06_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y06_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y06_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y06_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y06_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y06_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y06_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y06_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y06_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y06_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y06_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y06_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y06_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y06_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y06_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y06_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y06_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y06_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y06_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y06_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y06_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y06_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y06_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y06_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y06_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y06_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y06_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y06_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y06_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y06_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y06_SB_T4_WEST_SB_OUT_B16;
wire Tile_X03_Y06_clk_out;
wire [31:0] Tile_X03_Y06_config_out_config_addr;
wire [31:0] Tile_X03_Y06_config_out_config_data;
wire [0:0] Tile_X03_Y06_config_out_read;
wire [0:0] Tile_X03_Y06_config_out_write;
wire [8:0] Tile_X03_Y06_hi_unq1;
wire [7:0] Tile_X03_Y06_lo_unq1;
wire [31:0] Tile_X03_Y06_read_config_data;
wire Tile_X03_Y06_reset_out;
wire [0:0] Tile_X03_Y06_stall_out;
wire [8:0] Tile_X03_Y06_hi_out;
wire [7:0] Tile_X03_Y06_lo_out;
wire [15:0] Tile_X03_Y06_tile_id_in;
wire [0:0] Tile_X03_Y07_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y07_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y07_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y07_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y07_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y07_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y07_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y07_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y07_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y07_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y07_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y07_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y07_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y07_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y07_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y07_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y07_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y07_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y07_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y07_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y07_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y07_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y07_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y07_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y07_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y07_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y07_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y07_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y07_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y07_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y07_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y07_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y07_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y07_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y07_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y07_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y07_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y07_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y07_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y07_SB_T4_WEST_SB_OUT_B16;
wire Tile_X03_Y07_clk_out;
wire [31:0] Tile_X03_Y07_config_out_config_addr;
wire [31:0] Tile_X03_Y07_config_out_config_data;
wire [0:0] Tile_X03_Y07_config_out_read;
wire [0:0] Tile_X03_Y07_config_out_write;
wire [8:0] Tile_X03_Y07_hi_unq1;
wire [7:0] Tile_X03_Y07_lo_unq1;
wire [31:0] Tile_X03_Y07_read_config_data;
wire Tile_X03_Y07_reset_out;
wire [0:0] Tile_X03_Y07_stall_out;
wire [8:0] Tile_X03_Y07_hi_out;
wire [7:0] Tile_X03_Y07_lo_out;
wire [15:0] Tile_X03_Y07_tile_id_in;
wire [0:0] Tile_X03_Y08_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y08_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y08_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y08_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y08_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y08_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y08_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y08_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y08_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y08_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y08_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y08_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y08_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y08_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y08_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y08_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y08_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y08_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y08_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y08_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y08_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y08_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y08_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y08_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y08_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y08_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y08_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y08_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y08_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y08_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y08_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y08_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y08_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y08_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y08_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y08_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y08_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y08_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y08_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y08_SB_T4_WEST_SB_OUT_B16;
wire Tile_X03_Y08_clk_out;
wire [31:0] Tile_X03_Y08_config_out_config_addr;
wire [31:0] Tile_X03_Y08_config_out_config_data;
wire [0:0] Tile_X03_Y08_config_out_read;
wire [0:0] Tile_X03_Y08_config_out_write;
wire [8:0] Tile_X03_Y08_hi_unq1;
wire [7:0] Tile_X03_Y08_lo_unq1;
wire [31:0] Tile_X03_Y08_read_config_data;
wire Tile_X03_Y08_reset_out;
wire [0:0] Tile_X03_Y08_stall_out;
wire [8:0] Tile_X03_Y08_hi_out;
wire [7:0] Tile_X03_Y08_lo_out;
wire [15:0] Tile_X03_Y08_tile_id_in;
wire [0:0] Tile_X03_Y09_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y09_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y09_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y09_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y09_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y09_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y09_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y09_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y09_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y09_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y09_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y09_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y09_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y09_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y09_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y09_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y09_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y09_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y09_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y09_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y09_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y09_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y09_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y09_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y09_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y09_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y09_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y09_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y09_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y09_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y09_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y09_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y09_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y09_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y09_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y09_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y09_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y09_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y09_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y09_SB_T4_WEST_SB_OUT_B16;
wire Tile_X03_Y09_clk_out;
wire [31:0] Tile_X03_Y09_config_out_config_addr;
wire [31:0] Tile_X03_Y09_config_out_config_data;
wire [0:0] Tile_X03_Y09_config_out_read;
wire [0:0] Tile_X03_Y09_config_out_write;
wire [8:0] Tile_X03_Y09_hi_unq1;
wire [7:0] Tile_X03_Y09_lo_unq1;
wire [31:0] Tile_X03_Y09_read_config_data;
wire Tile_X03_Y09_reset_out;
wire [0:0] Tile_X03_Y09_stall_out;
wire [8:0] Tile_X03_Y09_hi_out;
wire [7:0] Tile_X03_Y09_lo_out;
wire [15:0] Tile_X03_Y09_tile_id_in;
wire [0:0] Tile_X03_Y0A_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0A_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0A_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0A_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0A_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0A_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0A_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0A_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0A_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0A_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0A_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0A_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0A_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0A_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0A_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0A_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0A_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0A_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0A_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0A_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0A_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0A_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0A_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0A_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0A_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0A_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0A_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0A_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0A_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0A_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0A_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0A_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0A_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0A_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0A_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0A_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0A_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0A_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0A_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0A_SB_T4_WEST_SB_OUT_B16;
wire Tile_X03_Y0A_clk_out;
wire [31:0] Tile_X03_Y0A_config_out_config_addr;
wire [31:0] Tile_X03_Y0A_config_out_config_data;
wire [0:0] Tile_X03_Y0A_config_out_read;
wire [0:0] Tile_X03_Y0A_config_out_write;
wire [8:0] Tile_X03_Y0A_hi_unq1;
wire [7:0] Tile_X03_Y0A_lo_unq1;
wire [31:0] Tile_X03_Y0A_read_config_data;
wire Tile_X03_Y0A_reset_out;
wire [0:0] Tile_X03_Y0A_stall_out;
wire [8:0] Tile_X03_Y0A_hi_out;
wire [7:0] Tile_X03_Y0A_lo_out;
wire [15:0] Tile_X03_Y0A_tile_id_in;
wire [0:0] Tile_X03_Y0B_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0B_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0B_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0B_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0B_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0B_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0B_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0B_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0B_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0B_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0B_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0B_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0B_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0B_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0B_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0B_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0B_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0B_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0B_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0B_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0B_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0B_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0B_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0B_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0B_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0B_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0B_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0B_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0B_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0B_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0B_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0B_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0B_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0B_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0B_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0B_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0B_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0B_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0B_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0B_SB_T4_WEST_SB_OUT_B16;
wire Tile_X03_Y0B_clk_out;
wire [31:0] Tile_X03_Y0B_config_out_config_addr;
wire [31:0] Tile_X03_Y0B_config_out_config_data;
wire [0:0] Tile_X03_Y0B_config_out_read;
wire [0:0] Tile_X03_Y0B_config_out_write;
wire [8:0] Tile_X03_Y0B_hi_unq1;
wire [7:0] Tile_X03_Y0B_lo_unq1;
wire [31:0] Tile_X03_Y0B_read_config_data;
wire Tile_X03_Y0B_reset_out;
wire [0:0] Tile_X03_Y0B_stall_out;
wire [8:0] Tile_X03_Y0B_hi_out;
wire [7:0] Tile_X03_Y0B_lo_out;
wire [15:0] Tile_X03_Y0B_tile_id_in;
wire [0:0] Tile_X03_Y0C_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0C_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0C_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0C_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0C_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0C_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0C_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0C_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0C_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0C_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0C_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0C_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0C_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0C_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0C_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0C_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0C_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0C_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0C_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0C_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0C_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0C_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0C_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0C_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0C_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0C_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0C_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0C_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0C_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0C_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0C_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0C_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0C_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0C_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0C_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0C_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0C_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0C_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0C_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0C_SB_T4_WEST_SB_OUT_B16;
wire Tile_X03_Y0C_clk_out;
wire [31:0] Tile_X03_Y0C_config_out_config_addr;
wire [31:0] Tile_X03_Y0C_config_out_config_data;
wire [0:0] Tile_X03_Y0C_config_out_read;
wire [0:0] Tile_X03_Y0C_config_out_write;
wire [8:0] Tile_X03_Y0C_hi_unq1;
wire [7:0] Tile_X03_Y0C_lo_unq1;
wire [31:0] Tile_X03_Y0C_read_config_data;
wire Tile_X03_Y0C_reset_out;
wire [0:0] Tile_X03_Y0C_stall_out;
wire [8:0] Tile_X03_Y0C_hi_out;
wire [7:0] Tile_X03_Y0C_lo_out;
wire [15:0] Tile_X03_Y0C_tile_id_in;
wire [0:0] Tile_X03_Y0D_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0D_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0D_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0D_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0D_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0D_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0D_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0D_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0D_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0D_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0D_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0D_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0D_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0D_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0D_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0D_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0D_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0D_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0D_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0D_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0D_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0D_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0D_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0D_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0D_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0D_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0D_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0D_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0D_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0D_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0D_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0D_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0D_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0D_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0D_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0D_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0D_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0D_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0D_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0D_SB_T4_WEST_SB_OUT_B16;
wire Tile_X03_Y0D_clk_out;
wire [31:0] Tile_X03_Y0D_config_out_config_addr;
wire [31:0] Tile_X03_Y0D_config_out_config_data;
wire [0:0] Tile_X03_Y0D_config_out_read;
wire [0:0] Tile_X03_Y0D_config_out_write;
wire [8:0] Tile_X03_Y0D_hi_unq1;
wire [7:0] Tile_X03_Y0D_lo_unq1;
wire [31:0] Tile_X03_Y0D_read_config_data;
wire Tile_X03_Y0D_reset_out;
wire [0:0] Tile_X03_Y0D_stall_out;
wire [8:0] Tile_X03_Y0D_hi_out;
wire [7:0] Tile_X03_Y0D_lo_out;
wire [15:0] Tile_X03_Y0D_tile_id_in;
wire [0:0] Tile_X03_Y0E_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0E_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0E_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0E_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0E_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0E_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0E_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0E_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0E_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0E_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0E_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0E_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0E_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0E_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0E_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0E_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0E_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0E_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0E_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0E_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0E_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0E_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0E_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0E_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0E_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0E_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0E_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0E_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0E_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0E_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0E_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0E_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0E_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0E_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0E_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0E_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0E_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0E_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0E_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0E_SB_T4_WEST_SB_OUT_B16;
wire Tile_X03_Y0E_clk_out;
wire [31:0] Tile_X03_Y0E_config_out_config_addr;
wire [31:0] Tile_X03_Y0E_config_out_config_data;
wire [0:0] Tile_X03_Y0E_config_out_read;
wire [0:0] Tile_X03_Y0E_config_out_write;
wire [8:0] Tile_X03_Y0E_hi_unq1;
wire [7:0] Tile_X03_Y0E_lo_unq1;
wire [31:0] Tile_X03_Y0E_read_config_data;
wire Tile_X03_Y0E_reset_out;
wire [0:0] Tile_X03_Y0E_stall_out;
wire [8:0] Tile_X03_Y0E_hi_out;
wire [7:0] Tile_X03_Y0E_lo_out;
wire [15:0] Tile_X03_Y0E_tile_id_in;
wire [0:0] Tile_X03_Y0F_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0F_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0F_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0F_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0F_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0F_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0F_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0F_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0F_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0F_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0F_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0F_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0F_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0F_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0F_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0F_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0F_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0F_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0F_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0F_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0F_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0F_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0F_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0F_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0F_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0F_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0F_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0F_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0F_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0F_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0F_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0F_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0F_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0F_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y0F_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0F_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0F_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y0F_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y0F_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y0F_SB_T4_WEST_SB_OUT_B16;
wire Tile_X03_Y0F_clk_out;
wire [31:0] Tile_X03_Y0F_config_out_config_addr;
wire [31:0] Tile_X03_Y0F_config_out_config_data;
wire [0:0] Tile_X03_Y0F_config_out_read;
wire [0:0] Tile_X03_Y0F_config_out_write;
wire [8:0] Tile_X03_Y0F_hi_unq1;
wire [7:0] Tile_X03_Y0F_lo_unq1;
wire [31:0] Tile_X03_Y0F_read_config_data;
wire Tile_X03_Y0F_reset_out;
wire [0:0] Tile_X03_Y0F_stall_out;
wire [8:0] Tile_X03_Y0F_hi_out;
wire [7:0] Tile_X03_Y0F_lo_out;
wire [15:0] Tile_X03_Y0F_tile_id_in;
wire [0:0] Tile_X03_Y10_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y10_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y10_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y10_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y10_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y10_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y10_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y10_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y10_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y10_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y10_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y10_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y10_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y10_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y10_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y10_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y10_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y10_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y10_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y10_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y10_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y10_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y10_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y10_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y10_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y10_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y10_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y10_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y10_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y10_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y10_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y10_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X03_Y10_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X03_Y10_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X03_Y10_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y10_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y10_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X03_Y10_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X03_Y10_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X03_Y10_SB_T4_WEST_SB_OUT_B16;
wire Tile_X03_Y10_clk_out;
wire [31:0] Tile_X03_Y10_config_out_config_addr;
wire [31:0] Tile_X03_Y10_config_out_config_data;
wire [0:0] Tile_X03_Y10_config_out_read;
wire [0:0] Tile_X03_Y10_config_out_write;
wire [8:0] Tile_X03_Y10_hi_unq1;
wire [7:0] Tile_X03_Y10_lo_unq1;
wire [31:0] Tile_X03_Y10_read_config_data;
wire Tile_X03_Y10_reset_out;
wire [0:0] Tile_X03_Y10_stall_out;
wire [8:0] Tile_X03_Y10_hi_out;
wire [7:0] Tile_X03_Y10_lo_out;
wire [15:0] Tile_X03_Y10_tile_id_in;
wire [0:0] Tile_X04_Y00_io2glb_1;
wire [0:0] Tile_X04_Y00_io2f_1;
wire [15:0] Tile_X04_Y00_io2glb_16;
wire [15:0] Tile_X04_Y00_io2f_16;
wire [8:0] Tile_X04_Y00_hi;
wire [7:0] Tile_X04_Y00_lo;
wire [0:0] Tile_X04_Y01_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y01_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y01_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y01_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y01_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y01_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y01_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y01_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y01_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y01_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y01_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y01_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y01_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y01_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y01_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y01_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y01_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y01_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y01_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y01_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y01_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y01_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y01_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y01_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y01_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y01_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y01_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y01_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y01_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y01_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y01_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y01_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y01_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y01_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y01_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y01_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y01_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y01_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y01_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y01_SB_T4_WEST_SB_OUT_B16;
wire Tile_X04_Y01_clk_out;
wire Tile_X04_Y01_clk_pass_through_out_bot;
wire Tile_X04_Y01_clk_pass_through_out_right;
wire [31:0] Tile_X04_Y01_config_out_config_addr;
wire [31:0] Tile_X04_Y01_config_out_config_data;
wire [0:0] Tile_X04_Y01_config_out_read;
wire [0:0] Tile_X04_Y01_config_out_write;
wire [8:0] Tile_X04_Y01_hi;
wire [7:0] Tile_X04_Y01_lo_unq1;
wire [31:0] Tile_X04_Y01_read_config_data;
wire Tile_X04_Y01_reset_out;
wire [0:0] Tile_X04_Y01_stall_out;
wire [7:0] Tile_X04_Y01_lo_out;
wire [15:0] Tile_X04_Y01_tile_id_in;
wire [0:0] Tile_X04_Y02_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y02_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y02_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y02_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y02_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y02_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y02_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y02_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y02_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y02_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y02_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y02_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y02_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y02_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y02_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y02_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y02_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y02_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y02_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y02_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y02_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y02_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y02_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y02_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y02_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y02_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y02_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y02_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y02_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y02_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y02_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y02_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y02_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y02_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y02_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y02_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y02_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y02_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y02_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y02_SB_T4_WEST_SB_OUT_B16;
wire Tile_X04_Y02_clk_out;
wire Tile_X04_Y02_clk_pass_through_out_bot;
wire Tile_X04_Y02_clk_pass_through_out_right;
wire [31:0] Tile_X04_Y02_config_out_config_addr;
wire [31:0] Tile_X04_Y02_config_out_config_data;
wire [0:0] Tile_X04_Y02_config_out_read;
wire [0:0] Tile_X04_Y02_config_out_write;
wire [8:0] Tile_X04_Y02_hi;
wire [7:0] Tile_X04_Y02_lo_unq1;
wire [31:0] Tile_X04_Y02_read_config_data;
wire Tile_X04_Y02_reset_out;
wire [0:0] Tile_X04_Y02_stall_out;
wire [7:0] Tile_X04_Y02_lo_out;
wire [15:0] Tile_X04_Y02_tile_id_in;
wire [0:0] Tile_X04_Y03_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y03_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y03_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y03_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y03_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y03_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y03_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y03_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y03_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y03_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y03_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y03_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y03_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y03_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y03_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y03_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y03_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y03_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y03_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y03_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y03_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y03_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y03_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y03_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y03_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y03_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y03_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y03_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y03_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y03_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y03_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y03_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y03_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y03_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y03_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y03_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y03_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y03_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y03_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y03_SB_T4_WEST_SB_OUT_B16;
wire Tile_X04_Y03_clk_out;
wire Tile_X04_Y03_clk_pass_through_out_bot;
wire Tile_X04_Y03_clk_pass_through_out_right;
wire [31:0] Tile_X04_Y03_config_out_config_addr;
wire [31:0] Tile_X04_Y03_config_out_config_data;
wire [0:0] Tile_X04_Y03_config_out_read;
wire [0:0] Tile_X04_Y03_config_out_write;
wire [8:0] Tile_X04_Y03_hi_unq1;
wire [7:0] Tile_X04_Y03_lo_unq1;
wire [31:0] Tile_X04_Y03_read_config_data;
wire Tile_X04_Y03_reset_out;
wire [0:0] Tile_X04_Y03_stall_out;
wire [8:0] Tile_X04_Y03_hi_out;
wire [7:0] Tile_X04_Y03_lo_out;
wire [15:0] Tile_X04_Y03_tile_id_in;
wire [0:0] Tile_X04_Y04_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y04_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y04_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y04_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y04_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y04_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y04_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y04_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y04_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y04_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y04_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y04_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y04_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y04_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y04_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y04_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y04_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y04_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y04_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y04_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y04_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y04_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y04_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y04_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y04_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y04_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y04_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y04_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y04_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y04_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y04_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y04_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y04_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y04_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y04_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y04_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y04_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y04_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y04_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y04_SB_T4_WEST_SB_OUT_B16;
wire Tile_X04_Y04_clk_out;
wire Tile_X04_Y04_clk_pass_through_out_bot;
wire Tile_X04_Y04_clk_pass_through_out_right;
wire [31:0] Tile_X04_Y04_config_out_config_addr;
wire [31:0] Tile_X04_Y04_config_out_config_data;
wire [0:0] Tile_X04_Y04_config_out_read;
wire [0:0] Tile_X04_Y04_config_out_write;
wire [8:0] Tile_X04_Y04_hi;
wire [7:0] Tile_X04_Y04_lo_unq1;
wire [31:0] Tile_X04_Y04_read_config_data;
wire Tile_X04_Y04_reset_out;
wire [0:0] Tile_X04_Y04_stall_out;
wire [7:0] Tile_X04_Y04_lo_out;
wire [15:0] Tile_X04_Y04_tile_id_in;
wire [0:0] Tile_X04_Y05_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y05_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y05_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y05_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y05_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y05_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y05_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y05_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y05_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y05_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y05_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y05_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y05_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y05_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y05_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y05_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y05_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y05_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y05_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y05_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y05_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y05_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y05_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y05_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y05_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y05_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y05_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y05_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y05_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y05_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y05_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y05_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y05_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y05_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y05_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y05_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y05_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y05_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y05_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y05_SB_T4_WEST_SB_OUT_B16;
wire Tile_X04_Y05_clk_out;
wire Tile_X04_Y05_clk_pass_through_out_bot;
wire Tile_X04_Y05_clk_pass_through_out_right;
wire [31:0] Tile_X04_Y05_config_out_config_addr;
wire [31:0] Tile_X04_Y05_config_out_config_data;
wire [0:0] Tile_X04_Y05_config_out_read;
wire [0:0] Tile_X04_Y05_config_out_write;
wire [8:0] Tile_X04_Y05_hi;
wire [7:0] Tile_X04_Y05_lo_unq1;
wire [31:0] Tile_X04_Y05_read_config_data;
wire Tile_X04_Y05_reset_out;
wire [0:0] Tile_X04_Y05_stall_out;
wire [7:0] Tile_X04_Y05_lo_out;
wire [15:0] Tile_X04_Y05_tile_id_in;
wire [0:0] Tile_X04_Y06_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y06_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y06_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y06_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y06_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y06_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y06_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y06_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y06_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y06_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y06_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y06_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y06_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y06_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y06_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y06_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y06_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y06_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y06_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y06_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y06_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y06_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y06_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y06_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y06_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y06_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y06_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y06_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y06_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y06_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y06_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y06_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y06_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y06_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y06_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y06_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y06_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y06_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y06_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y06_SB_T4_WEST_SB_OUT_B16;
wire Tile_X04_Y06_clk_out;
wire Tile_X04_Y06_clk_pass_through_out_bot;
wire Tile_X04_Y06_clk_pass_through_out_right;
wire [31:0] Tile_X04_Y06_config_out_config_addr;
wire [31:0] Tile_X04_Y06_config_out_config_data;
wire [0:0] Tile_X04_Y06_config_out_read;
wire [0:0] Tile_X04_Y06_config_out_write;
wire [8:0] Tile_X04_Y06_hi;
wire [7:0] Tile_X04_Y06_lo_unq1;
wire [31:0] Tile_X04_Y06_read_config_data;
wire Tile_X04_Y06_reset_out;
wire [0:0] Tile_X04_Y06_stall_out;
wire [7:0] Tile_X04_Y06_lo_out;
wire [15:0] Tile_X04_Y06_tile_id_in;
wire [0:0] Tile_X04_Y07_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y07_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y07_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y07_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y07_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y07_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y07_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y07_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y07_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y07_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y07_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y07_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y07_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y07_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y07_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y07_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y07_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y07_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y07_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y07_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y07_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y07_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y07_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y07_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y07_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y07_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y07_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y07_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y07_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y07_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y07_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y07_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y07_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y07_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y07_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y07_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y07_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y07_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y07_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y07_SB_T4_WEST_SB_OUT_B16;
wire Tile_X04_Y07_clk_out;
wire Tile_X04_Y07_clk_pass_through_out_bot;
wire Tile_X04_Y07_clk_pass_through_out_right;
wire [31:0] Tile_X04_Y07_config_out_config_addr;
wire [31:0] Tile_X04_Y07_config_out_config_data;
wire [0:0] Tile_X04_Y07_config_out_read;
wire [0:0] Tile_X04_Y07_config_out_write;
wire [8:0] Tile_X04_Y07_hi_unq1;
wire [7:0] Tile_X04_Y07_lo_unq1;
wire [31:0] Tile_X04_Y07_read_config_data;
wire Tile_X04_Y07_reset_out;
wire [0:0] Tile_X04_Y07_stall_out;
wire [8:0] Tile_X04_Y07_hi_out;
wire [7:0] Tile_X04_Y07_lo_out;
wire [15:0] Tile_X04_Y07_tile_id_in;
wire [0:0] Tile_X04_Y08_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y08_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y08_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y08_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y08_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y08_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y08_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y08_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y08_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y08_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y08_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y08_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y08_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y08_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y08_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y08_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y08_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y08_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y08_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y08_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y08_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y08_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y08_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y08_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y08_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y08_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y08_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y08_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y08_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y08_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y08_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y08_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y08_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y08_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y08_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y08_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y08_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y08_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y08_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y08_SB_T4_WEST_SB_OUT_B16;
wire Tile_X04_Y08_clk_out;
wire Tile_X04_Y08_clk_pass_through_out_bot;
wire Tile_X04_Y08_clk_pass_through_out_right;
wire [31:0] Tile_X04_Y08_config_out_config_addr;
wire [31:0] Tile_X04_Y08_config_out_config_data;
wire [0:0] Tile_X04_Y08_config_out_read;
wire [0:0] Tile_X04_Y08_config_out_write;
wire [8:0] Tile_X04_Y08_hi;
wire [7:0] Tile_X04_Y08_lo_unq1;
wire [31:0] Tile_X04_Y08_read_config_data;
wire Tile_X04_Y08_reset_out;
wire [0:0] Tile_X04_Y08_stall_out;
wire [7:0] Tile_X04_Y08_lo_out;
wire [15:0] Tile_X04_Y08_tile_id_in;
wire [0:0] Tile_X04_Y09_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y09_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y09_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y09_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y09_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y09_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y09_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y09_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y09_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y09_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y09_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y09_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y09_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y09_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y09_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y09_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y09_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y09_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y09_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y09_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y09_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y09_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y09_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y09_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y09_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y09_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y09_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y09_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y09_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y09_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y09_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y09_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y09_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y09_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y09_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y09_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y09_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y09_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y09_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y09_SB_T4_WEST_SB_OUT_B16;
wire Tile_X04_Y09_clk_out;
wire Tile_X04_Y09_clk_pass_through_out_bot;
wire Tile_X04_Y09_clk_pass_through_out_right;
wire [31:0] Tile_X04_Y09_config_out_config_addr;
wire [31:0] Tile_X04_Y09_config_out_config_data;
wire [0:0] Tile_X04_Y09_config_out_read;
wire [0:0] Tile_X04_Y09_config_out_write;
wire [8:0] Tile_X04_Y09_hi;
wire [7:0] Tile_X04_Y09_lo_unq1;
wire [31:0] Tile_X04_Y09_read_config_data;
wire Tile_X04_Y09_reset_out;
wire [0:0] Tile_X04_Y09_stall_out;
wire [7:0] Tile_X04_Y09_lo_out;
wire [15:0] Tile_X04_Y09_tile_id_in;
wire [0:0] Tile_X04_Y0A_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0A_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0A_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0A_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0A_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0A_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0A_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0A_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0A_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0A_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0A_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0A_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0A_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0A_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0A_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0A_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0A_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0A_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0A_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0A_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0A_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0A_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0A_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0A_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0A_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0A_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0A_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0A_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0A_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0A_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0A_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0A_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0A_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0A_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0A_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0A_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0A_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0A_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0A_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0A_SB_T4_WEST_SB_OUT_B16;
wire Tile_X04_Y0A_clk_out;
wire Tile_X04_Y0A_clk_pass_through_out_bot;
wire Tile_X04_Y0A_clk_pass_through_out_right;
wire [31:0] Tile_X04_Y0A_config_out_config_addr;
wire [31:0] Tile_X04_Y0A_config_out_config_data;
wire [0:0] Tile_X04_Y0A_config_out_read;
wire [0:0] Tile_X04_Y0A_config_out_write;
wire [8:0] Tile_X04_Y0A_hi;
wire [7:0] Tile_X04_Y0A_lo_unq1;
wire [31:0] Tile_X04_Y0A_read_config_data;
wire Tile_X04_Y0A_reset_out;
wire [0:0] Tile_X04_Y0A_stall_out;
wire [7:0] Tile_X04_Y0A_lo_out;
wire [15:0] Tile_X04_Y0A_tile_id_in;
wire [0:0] Tile_X04_Y0B_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0B_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0B_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0B_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0B_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0B_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0B_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0B_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0B_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0B_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0B_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0B_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0B_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0B_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0B_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0B_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0B_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0B_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0B_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0B_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0B_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0B_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0B_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0B_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0B_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0B_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0B_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0B_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0B_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0B_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0B_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0B_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0B_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0B_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0B_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0B_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0B_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0B_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0B_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0B_SB_T4_WEST_SB_OUT_B16;
wire Tile_X04_Y0B_clk_out;
wire Tile_X04_Y0B_clk_pass_through_out_bot;
wire Tile_X04_Y0B_clk_pass_through_out_right;
wire [31:0] Tile_X04_Y0B_config_out_config_addr;
wire [31:0] Tile_X04_Y0B_config_out_config_data;
wire [0:0] Tile_X04_Y0B_config_out_read;
wire [0:0] Tile_X04_Y0B_config_out_write;
wire [8:0] Tile_X04_Y0B_hi_unq1;
wire [7:0] Tile_X04_Y0B_lo_unq1;
wire [31:0] Tile_X04_Y0B_read_config_data;
wire Tile_X04_Y0B_reset_out;
wire [0:0] Tile_X04_Y0B_stall_out;
wire [8:0] Tile_X04_Y0B_hi_out;
wire [7:0] Tile_X04_Y0B_lo_out;
wire [15:0] Tile_X04_Y0B_tile_id_in;
wire [0:0] Tile_X04_Y0C_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0C_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0C_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0C_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0C_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0C_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0C_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0C_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0C_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0C_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0C_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0C_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0C_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0C_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0C_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0C_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0C_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0C_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0C_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0C_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0C_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0C_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0C_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0C_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0C_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0C_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0C_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0C_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0C_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0C_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0C_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0C_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0C_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0C_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0C_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0C_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0C_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0C_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0C_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0C_SB_T4_WEST_SB_OUT_B16;
wire Tile_X04_Y0C_clk_out;
wire Tile_X04_Y0C_clk_pass_through_out_bot;
wire Tile_X04_Y0C_clk_pass_through_out_right;
wire [31:0] Tile_X04_Y0C_config_out_config_addr;
wire [31:0] Tile_X04_Y0C_config_out_config_data;
wire [0:0] Tile_X04_Y0C_config_out_read;
wire [0:0] Tile_X04_Y0C_config_out_write;
wire [8:0] Tile_X04_Y0C_hi_unq1;
wire [7:0] Tile_X04_Y0C_lo_unq1;
wire [31:0] Tile_X04_Y0C_read_config_data;
wire Tile_X04_Y0C_reset_out;
wire [0:0] Tile_X04_Y0C_stall_out;
wire [8:0] Tile_X04_Y0C_hi_out;
wire [7:0] Tile_X04_Y0C_lo_out;
wire [15:0] Tile_X04_Y0C_tile_id_in;
wire [0:0] Tile_X04_Y0D_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0D_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0D_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0D_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0D_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0D_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0D_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0D_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0D_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0D_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0D_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0D_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0D_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0D_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0D_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0D_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0D_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0D_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0D_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0D_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0D_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0D_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0D_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0D_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0D_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0D_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0D_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0D_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0D_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0D_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0D_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0D_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0D_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0D_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0D_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0D_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0D_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0D_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0D_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0D_SB_T4_WEST_SB_OUT_B16;
wire Tile_X04_Y0D_clk_out;
wire Tile_X04_Y0D_clk_pass_through_out_bot;
wire Tile_X04_Y0D_clk_pass_through_out_right;
wire [31:0] Tile_X04_Y0D_config_out_config_addr;
wire [31:0] Tile_X04_Y0D_config_out_config_data;
wire [0:0] Tile_X04_Y0D_config_out_read;
wire [0:0] Tile_X04_Y0D_config_out_write;
wire [8:0] Tile_X04_Y0D_hi_unq1;
wire [7:0] Tile_X04_Y0D_lo_unq1;
wire [31:0] Tile_X04_Y0D_read_config_data;
wire Tile_X04_Y0D_reset_out;
wire [0:0] Tile_X04_Y0D_stall_out;
wire [8:0] Tile_X04_Y0D_hi_out;
wire [7:0] Tile_X04_Y0D_lo_out;
wire [15:0] Tile_X04_Y0D_tile_id_in;
wire [0:0] Tile_X04_Y0E_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0E_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0E_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0E_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0E_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0E_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0E_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0E_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0E_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0E_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0E_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0E_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0E_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0E_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0E_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0E_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0E_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0E_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0E_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0E_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0E_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0E_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0E_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0E_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0E_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0E_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0E_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0E_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0E_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0E_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0E_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0E_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0E_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0E_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0E_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0E_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0E_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0E_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0E_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0E_SB_T4_WEST_SB_OUT_B16;
wire Tile_X04_Y0E_clk_out;
wire Tile_X04_Y0E_clk_pass_through_out_bot;
wire Tile_X04_Y0E_clk_pass_through_out_right;
wire [31:0] Tile_X04_Y0E_config_out_config_addr;
wire [31:0] Tile_X04_Y0E_config_out_config_data;
wire [0:0] Tile_X04_Y0E_config_out_read;
wire [0:0] Tile_X04_Y0E_config_out_write;
wire [8:0] Tile_X04_Y0E_hi_unq1;
wire [7:0] Tile_X04_Y0E_lo_unq1;
wire [31:0] Tile_X04_Y0E_read_config_data;
wire Tile_X04_Y0E_reset_out;
wire [0:0] Tile_X04_Y0E_stall_out;
wire [8:0] Tile_X04_Y0E_hi_out;
wire [7:0] Tile_X04_Y0E_lo_out;
wire [15:0] Tile_X04_Y0E_tile_id_in;
wire [0:0] Tile_X04_Y0F_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0F_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0F_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0F_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0F_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0F_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0F_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0F_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0F_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0F_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0F_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0F_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0F_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0F_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0F_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0F_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0F_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0F_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0F_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0F_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0F_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0F_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0F_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0F_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0F_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0F_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0F_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0F_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0F_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0F_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0F_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0F_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0F_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0F_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y0F_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0F_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0F_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y0F_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y0F_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y0F_SB_T4_WEST_SB_OUT_B16;
wire Tile_X04_Y0F_clk_out;
wire Tile_X04_Y0F_clk_pass_through_out_bot;
wire Tile_X04_Y0F_clk_pass_through_out_right;
wire [31:0] Tile_X04_Y0F_config_out_config_addr;
wire [31:0] Tile_X04_Y0F_config_out_config_data;
wire [0:0] Tile_X04_Y0F_config_out_read;
wire [0:0] Tile_X04_Y0F_config_out_write;
wire [8:0] Tile_X04_Y0F_hi_unq1;
wire [7:0] Tile_X04_Y0F_lo_unq1;
wire [31:0] Tile_X04_Y0F_read_config_data;
wire Tile_X04_Y0F_reset_out;
wire [0:0] Tile_X04_Y0F_stall_out;
wire [8:0] Tile_X04_Y0F_hi_out;
wire [7:0] Tile_X04_Y0F_lo_out;
wire [15:0] Tile_X04_Y0F_tile_id_in;
wire [0:0] Tile_X04_Y10_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y10_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y10_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y10_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y10_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y10_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y10_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y10_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y10_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y10_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y10_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y10_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y10_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y10_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y10_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y10_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y10_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y10_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y10_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y10_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y10_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y10_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y10_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y10_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y10_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y10_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y10_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y10_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y10_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y10_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y10_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y10_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X04_Y10_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X04_Y10_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X04_Y10_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y10_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y10_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X04_Y10_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X04_Y10_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X04_Y10_SB_T4_WEST_SB_OUT_B16;
wire Tile_X04_Y10_clk_out;
wire Tile_X04_Y10_clk_pass_through_out_bot;
wire Tile_X04_Y10_clk_pass_through_out_right;
wire [31:0] Tile_X04_Y10_config_out_config_addr;
wire [31:0] Tile_X04_Y10_config_out_config_data;
wire [0:0] Tile_X04_Y10_config_out_read;
wire [0:0] Tile_X04_Y10_config_out_write;
wire [8:0] Tile_X04_Y10_hi;
wire [7:0] Tile_X04_Y10_lo_unq1;
wire [31:0] Tile_X04_Y10_read_config_data;
wire Tile_X04_Y10_reset_out;
wire [0:0] Tile_X04_Y10_stall_out;
wire [7:0] Tile_X04_Y10_lo_out;
wire [15:0] Tile_X04_Y10_tile_id_in;
wire [0:0] Tile_X05_Y00_io2glb_1;
wire [0:0] Tile_X05_Y00_io2f_1;
wire [15:0] Tile_X05_Y00_io2glb_16;
wire [15:0] Tile_X05_Y00_io2f_16;
wire [8:0] Tile_X05_Y00_hi;
wire [7:0] Tile_X05_Y00_lo;
wire [0:0] Tile_X05_Y01_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y01_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y01_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y01_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y01_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y01_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y01_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y01_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y01_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y01_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y01_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y01_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y01_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y01_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y01_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y01_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y01_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y01_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y01_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y01_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y01_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y01_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y01_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y01_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y01_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y01_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y01_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y01_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y01_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y01_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y01_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y01_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y01_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y01_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y01_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y01_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y01_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y01_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y01_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y01_SB_T4_WEST_SB_OUT_B16;
wire Tile_X05_Y01_clk_out;
wire Tile_X05_Y01_clk_pass_through_out_bot;
wire Tile_X05_Y01_clk_pass_through_out_right;
wire [31:0] Tile_X05_Y01_config_out_config_addr;
wire [31:0] Tile_X05_Y01_config_out_config_data;
wire [0:0] Tile_X05_Y01_config_out_read;
wire [0:0] Tile_X05_Y01_config_out_write;
wire [8:0] Tile_X05_Y01_hi;
wire [7:0] Tile_X05_Y01_lo_unq1;
wire [31:0] Tile_X05_Y01_read_config_data;
wire Tile_X05_Y01_reset_out;
wire [0:0] Tile_X05_Y01_stall_out;
wire [7:0] Tile_X05_Y01_lo_out;
wire [15:0] Tile_X05_Y01_tile_id_in;
wire [0:0] Tile_X05_Y02_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y02_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y02_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y02_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y02_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y02_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y02_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y02_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y02_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y02_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y02_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y02_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y02_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y02_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y02_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y02_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y02_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y02_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y02_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y02_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y02_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y02_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y02_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y02_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y02_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y02_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y02_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y02_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y02_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y02_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y02_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y02_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y02_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y02_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y02_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y02_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y02_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y02_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y02_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y02_SB_T4_WEST_SB_OUT_B16;
wire Tile_X05_Y02_clk_out;
wire Tile_X05_Y02_clk_pass_through_out_bot;
wire Tile_X05_Y02_clk_pass_through_out_right;
wire [31:0] Tile_X05_Y02_config_out_config_addr;
wire [31:0] Tile_X05_Y02_config_out_config_data;
wire [0:0] Tile_X05_Y02_config_out_read;
wire [0:0] Tile_X05_Y02_config_out_write;
wire [8:0] Tile_X05_Y02_hi;
wire [7:0] Tile_X05_Y02_lo_unq1;
wire [31:0] Tile_X05_Y02_read_config_data;
wire Tile_X05_Y02_reset_out;
wire [0:0] Tile_X05_Y02_stall_out;
wire [7:0] Tile_X05_Y02_lo_out;
wire [15:0] Tile_X05_Y02_tile_id_in;
wire [0:0] Tile_X05_Y03_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y03_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y03_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y03_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y03_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y03_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y03_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y03_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y03_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y03_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y03_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y03_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y03_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y03_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y03_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y03_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y03_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y03_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y03_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y03_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y03_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y03_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y03_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y03_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y03_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y03_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y03_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y03_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y03_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y03_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y03_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y03_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y03_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y03_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y03_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y03_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y03_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y03_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y03_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y03_SB_T4_WEST_SB_OUT_B16;
wire Tile_X05_Y03_clk_out;
wire Tile_X05_Y03_clk_pass_through_out_bot;
wire Tile_X05_Y03_clk_pass_through_out_right;
wire [31:0] Tile_X05_Y03_config_out_config_addr;
wire [31:0] Tile_X05_Y03_config_out_config_data;
wire [0:0] Tile_X05_Y03_config_out_read;
wire [0:0] Tile_X05_Y03_config_out_write;
wire [8:0] Tile_X05_Y03_hi_unq1;
wire [7:0] Tile_X05_Y03_lo_unq1;
wire [31:0] Tile_X05_Y03_read_config_data;
wire Tile_X05_Y03_reset_out;
wire [0:0] Tile_X05_Y03_stall_out;
wire [8:0] Tile_X05_Y03_hi_out;
wire [7:0] Tile_X05_Y03_lo_out;
wire [15:0] Tile_X05_Y03_tile_id_in;
wire [0:0] Tile_X05_Y04_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y04_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y04_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y04_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y04_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y04_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y04_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y04_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y04_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y04_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y04_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y04_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y04_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y04_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y04_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y04_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y04_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y04_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y04_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y04_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y04_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y04_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y04_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y04_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y04_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y04_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y04_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y04_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y04_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y04_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y04_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y04_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y04_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y04_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y04_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y04_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y04_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y04_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y04_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y04_SB_T4_WEST_SB_OUT_B16;
wire Tile_X05_Y04_clk_out;
wire Tile_X05_Y04_clk_pass_through_out_bot;
wire Tile_X05_Y04_clk_pass_through_out_right;
wire [31:0] Tile_X05_Y04_config_out_config_addr;
wire [31:0] Tile_X05_Y04_config_out_config_data;
wire [0:0] Tile_X05_Y04_config_out_read;
wire [0:0] Tile_X05_Y04_config_out_write;
wire [8:0] Tile_X05_Y04_hi;
wire [7:0] Tile_X05_Y04_lo_unq1;
wire [31:0] Tile_X05_Y04_read_config_data;
wire Tile_X05_Y04_reset_out;
wire [0:0] Tile_X05_Y04_stall_out;
wire [7:0] Tile_X05_Y04_lo_out;
wire [15:0] Tile_X05_Y04_tile_id_in;
wire [0:0] Tile_X05_Y05_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y05_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y05_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y05_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y05_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y05_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y05_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y05_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y05_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y05_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y05_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y05_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y05_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y05_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y05_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y05_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y05_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y05_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y05_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y05_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y05_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y05_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y05_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y05_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y05_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y05_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y05_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y05_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y05_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y05_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y05_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y05_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y05_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y05_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y05_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y05_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y05_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y05_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y05_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y05_SB_T4_WEST_SB_OUT_B16;
wire Tile_X05_Y05_clk_out;
wire Tile_X05_Y05_clk_pass_through_out_bot;
wire Tile_X05_Y05_clk_pass_through_out_right;
wire [31:0] Tile_X05_Y05_config_out_config_addr;
wire [31:0] Tile_X05_Y05_config_out_config_data;
wire [0:0] Tile_X05_Y05_config_out_read;
wire [0:0] Tile_X05_Y05_config_out_write;
wire [8:0] Tile_X05_Y05_hi;
wire [7:0] Tile_X05_Y05_lo_unq1;
wire [31:0] Tile_X05_Y05_read_config_data;
wire Tile_X05_Y05_reset_out;
wire [0:0] Tile_X05_Y05_stall_out;
wire [7:0] Tile_X05_Y05_lo_out;
wire [15:0] Tile_X05_Y05_tile_id_in;
wire [0:0] Tile_X05_Y06_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y06_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y06_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y06_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y06_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y06_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y06_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y06_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y06_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y06_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y06_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y06_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y06_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y06_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y06_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y06_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y06_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y06_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y06_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y06_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y06_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y06_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y06_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y06_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y06_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y06_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y06_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y06_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y06_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y06_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y06_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y06_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y06_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y06_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y06_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y06_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y06_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y06_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y06_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y06_SB_T4_WEST_SB_OUT_B16;
wire Tile_X05_Y06_clk_out;
wire Tile_X05_Y06_clk_pass_through_out_bot;
wire Tile_X05_Y06_clk_pass_through_out_right;
wire [31:0] Tile_X05_Y06_config_out_config_addr;
wire [31:0] Tile_X05_Y06_config_out_config_data;
wire [0:0] Tile_X05_Y06_config_out_read;
wire [0:0] Tile_X05_Y06_config_out_write;
wire [8:0] Tile_X05_Y06_hi;
wire [7:0] Tile_X05_Y06_lo_unq1;
wire [31:0] Tile_X05_Y06_read_config_data;
wire Tile_X05_Y06_reset_out;
wire [0:0] Tile_X05_Y06_stall_out;
wire [7:0] Tile_X05_Y06_lo_out;
wire [15:0] Tile_X05_Y06_tile_id_in;
wire [0:0] Tile_X05_Y07_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y07_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y07_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y07_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y07_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y07_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y07_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y07_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y07_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y07_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y07_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y07_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y07_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y07_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y07_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y07_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y07_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y07_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y07_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y07_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y07_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y07_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y07_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y07_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y07_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y07_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y07_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y07_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y07_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y07_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y07_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y07_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y07_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y07_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y07_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y07_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y07_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y07_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y07_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y07_SB_T4_WEST_SB_OUT_B16;
wire Tile_X05_Y07_clk_out;
wire Tile_X05_Y07_clk_pass_through_out_bot;
wire Tile_X05_Y07_clk_pass_through_out_right;
wire [31:0] Tile_X05_Y07_config_out_config_addr;
wire [31:0] Tile_X05_Y07_config_out_config_data;
wire [0:0] Tile_X05_Y07_config_out_read;
wire [0:0] Tile_X05_Y07_config_out_write;
wire [8:0] Tile_X05_Y07_hi_unq1;
wire [7:0] Tile_X05_Y07_lo_unq1;
wire [31:0] Tile_X05_Y07_read_config_data;
wire Tile_X05_Y07_reset_out;
wire [0:0] Tile_X05_Y07_stall_out;
wire [8:0] Tile_X05_Y07_hi_out;
wire [7:0] Tile_X05_Y07_lo_out;
wire [15:0] Tile_X05_Y07_tile_id_in;
wire [0:0] Tile_X05_Y08_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y08_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y08_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y08_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y08_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y08_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y08_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y08_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y08_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y08_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y08_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y08_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y08_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y08_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y08_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y08_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y08_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y08_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y08_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y08_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y08_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y08_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y08_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y08_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y08_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y08_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y08_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y08_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y08_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y08_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y08_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y08_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y08_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y08_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y08_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y08_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y08_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y08_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y08_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y08_SB_T4_WEST_SB_OUT_B16;
wire Tile_X05_Y08_clk_out;
wire Tile_X05_Y08_clk_pass_through_out_bot;
wire Tile_X05_Y08_clk_pass_through_out_right;
wire [31:0] Tile_X05_Y08_config_out_config_addr;
wire [31:0] Tile_X05_Y08_config_out_config_data;
wire [0:0] Tile_X05_Y08_config_out_read;
wire [0:0] Tile_X05_Y08_config_out_write;
wire [8:0] Tile_X05_Y08_hi;
wire [7:0] Tile_X05_Y08_lo_unq1;
wire [31:0] Tile_X05_Y08_read_config_data;
wire Tile_X05_Y08_reset_out;
wire [0:0] Tile_X05_Y08_stall_out;
wire [7:0] Tile_X05_Y08_lo_out;
wire [15:0] Tile_X05_Y08_tile_id_in;
wire [0:0] Tile_X05_Y09_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y09_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y09_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y09_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y09_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y09_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y09_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y09_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y09_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y09_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y09_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y09_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y09_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y09_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y09_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y09_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y09_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y09_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y09_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y09_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y09_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y09_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y09_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y09_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y09_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y09_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y09_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y09_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y09_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y09_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y09_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y09_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y09_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y09_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y09_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y09_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y09_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y09_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y09_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y09_SB_T4_WEST_SB_OUT_B16;
wire Tile_X05_Y09_clk_out;
wire Tile_X05_Y09_clk_pass_through_out_bot;
wire Tile_X05_Y09_clk_pass_through_out_right;
wire [31:0] Tile_X05_Y09_config_out_config_addr;
wire [31:0] Tile_X05_Y09_config_out_config_data;
wire [0:0] Tile_X05_Y09_config_out_read;
wire [0:0] Tile_X05_Y09_config_out_write;
wire [8:0] Tile_X05_Y09_hi;
wire [7:0] Tile_X05_Y09_lo_unq1;
wire [31:0] Tile_X05_Y09_read_config_data;
wire Tile_X05_Y09_reset_out;
wire [0:0] Tile_X05_Y09_stall_out;
wire [7:0] Tile_X05_Y09_lo_out;
wire [15:0] Tile_X05_Y09_tile_id_in;
wire [0:0] Tile_X05_Y0A_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0A_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0A_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0A_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0A_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0A_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0A_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0A_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0A_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0A_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0A_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0A_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0A_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0A_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0A_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0A_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0A_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0A_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0A_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0A_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0A_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0A_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0A_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0A_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0A_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0A_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0A_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0A_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0A_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0A_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0A_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0A_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0A_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0A_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0A_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0A_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0A_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0A_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0A_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0A_SB_T4_WEST_SB_OUT_B16;
wire Tile_X05_Y0A_clk_out;
wire Tile_X05_Y0A_clk_pass_through_out_bot;
wire Tile_X05_Y0A_clk_pass_through_out_right;
wire [31:0] Tile_X05_Y0A_config_out_config_addr;
wire [31:0] Tile_X05_Y0A_config_out_config_data;
wire [0:0] Tile_X05_Y0A_config_out_read;
wire [0:0] Tile_X05_Y0A_config_out_write;
wire [8:0] Tile_X05_Y0A_hi;
wire [7:0] Tile_X05_Y0A_lo_unq1;
wire [31:0] Tile_X05_Y0A_read_config_data;
wire Tile_X05_Y0A_reset_out;
wire [0:0] Tile_X05_Y0A_stall_out;
wire [7:0] Tile_X05_Y0A_lo_out;
wire [15:0] Tile_X05_Y0A_tile_id_in;
wire [0:0] Tile_X05_Y0B_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0B_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0B_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0B_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0B_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0B_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0B_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0B_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0B_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0B_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0B_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0B_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0B_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0B_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0B_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0B_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0B_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0B_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0B_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0B_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0B_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0B_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0B_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0B_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0B_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0B_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0B_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0B_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0B_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0B_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0B_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0B_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0B_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0B_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0B_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0B_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0B_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0B_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0B_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0B_SB_T4_WEST_SB_OUT_B16;
wire Tile_X05_Y0B_clk_out;
wire Tile_X05_Y0B_clk_pass_through_out_bot;
wire Tile_X05_Y0B_clk_pass_through_out_right;
wire [31:0] Tile_X05_Y0B_config_out_config_addr;
wire [31:0] Tile_X05_Y0B_config_out_config_data;
wire [0:0] Tile_X05_Y0B_config_out_read;
wire [0:0] Tile_X05_Y0B_config_out_write;
wire [8:0] Tile_X05_Y0B_hi_unq1;
wire [7:0] Tile_X05_Y0B_lo_unq1;
wire [31:0] Tile_X05_Y0B_read_config_data;
wire Tile_X05_Y0B_reset_out;
wire [0:0] Tile_X05_Y0B_stall_out;
wire [8:0] Tile_X05_Y0B_hi_out;
wire [7:0] Tile_X05_Y0B_lo_out;
wire [15:0] Tile_X05_Y0B_tile_id_in;
wire [0:0] Tile_X05_Y0C_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0C_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0C_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0C_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0C_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0C_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0C_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0C_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0C_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0C_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0C_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0C_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0C_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0C_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0C_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0C_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0C_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0C_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0C_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0C_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0C_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0C_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0C_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0C_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0C_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0C_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0C_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0C_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0C_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0C_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0C_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0C_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0C_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0C_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0C_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0C_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0C_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0C_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0C_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0C_SB_T4_WEST_SB_OUT_B16;
wire Tile_X05_Y0C_clk_out;
wire Tile_X05_Y0C_clk_pass_through_out_bot;
wire Tile_X05_Y0C_clk_pass_through_out_right;
wire [31:0] Tile_X05_Y0C_config_out_config_addr;
wire [31:0] Tile_X05_Y0C_config_out_config_data;
wire [0:0] Tile_X05_Y0C_config_out_read;
wire [0:0] Tile_X05_Y0C_config_out_write;
wire [8:0] Tile_X05_Y0C_hi_unq1;
wire [7:0] Tile_X05_Y0C_lo_unq1;
wire [31:0] Tile_X05_Y0C_read_config_data;
wire Tile_X05_Y0C_reset_out;
wire [0:0] Tile_X05_Y0C_stall_out;
wire [8:0] Tile_X05_Y0C_hi_out;
wire [7:0] Tile_X05_Y0C_lo_out;
wire [15:0] Tile_X05_Y0C_tile_id_in;
wire [0:0] Tile_X05_Y0D_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0D_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0D_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0D_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0D_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0D_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0D_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0D_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0D_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0D_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0D_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0D_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0D_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0D_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0D_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0D_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0D_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0D_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0D_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0D_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0D_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0D_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0D_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0D_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0D_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0D_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0D_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0D_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0D_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0D_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0D_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0D_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0D_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0D_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0D_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0D_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0D_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0D_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0D_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0D_SB_T4_WEST_SB_OUT_B16;
wire Tile_X05_Y0D_clk_out;
wire Tile_X05_Y0D_clk_pass_through_out_bot;
wire Tile_X05_Y0D_clk_pass_through_out_right;
wire [31:0] Tile_X05_Y0D_config_out_config_addr;
wire [31:0] Tile_X05_Y0D_config_out_config_data;
wire [0:0] Tile_X05_Y0D_config_out_read;
wire [0:0] Tile_X05_Y0D_config_out_write;
wire [8:0] Tile_X05_Y0D_hi_unq1;
wire [7:0] Tile_X05_Y0D_lo_unq1;
wire [31:0] Tile_X05_Y0D_read_config_data;
wire Tile_X05_Y0D_reset_out;
wire [0:0] Tile_X05_Y0D_stall_out;
wire [8:0] Tile_X05_Y0D_hi_out;
wire [7:0] Tile_X05_Y0D_lo_out;
wire [15:0] Tile_X05_Y0D_tile_id_in;
wire [0:0] Tile_X05_Y0E_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0E_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0E_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0E_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0E_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0E_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0E_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0E_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0E_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0E_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0E_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0E_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0E_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0E_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0E_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0E_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0E_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0E_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0E_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0E_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0E_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0E_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0E_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0E_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0E_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0E_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0E_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0E_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0E_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0E_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0E_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0E_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0E_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0E_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0E_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0E_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0E_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0E_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0E_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0E_SB_T4_WEST_SB_OUT_B16;
wire Tile_X05_Y0E_clk_out;
wire Tile_X05_Y0E_clk_pass_through_out_bot;
wire Tile_X05_Y0E_clk_pass_through_out_right;
wire [31:0] Tile_X05_Y0E_config_out_config_addr;
wire [31:0] Tile_X05_Y0E_config_out_config_data;
wire [0:0] Tile_X05_Y0E_config_out_read;
wire [0:0] Tile_X05_Y0E_config_out_write;
wire [8:0] Tile_X05_Y0E_hi_unq1;
wire [7:0] Tile_X05_Y0E_lo_unq1;
wire [31:0] Tile_X05_Y0E_read_config_data;
wire Tile_X05_Y0E_reset_out;
wire [0:0] Tile_X05_Y0E_stall_out;
wire [8:0] Tile_X05_Y0E_hi_out;
wire [7:0] Tile_X05_Y0E_lo_out;
wire [15:0] Tile_X05_Y0E_tile_id_in;
wire [0:0] Tile_X05_Y0F_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0F_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0F_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0F_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0F_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0F_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0F_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0F_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0F_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0F_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0F_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0F_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0F_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0F_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0F_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0F_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0F_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0F_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0F_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0F_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0F_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0F_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0F_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0F_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0F_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0F_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0F_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0F_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0F_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0F_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0F_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0F_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0F_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0F_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y0F_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0F_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0F_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y0F_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y0F_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y0F_SB_T4_WEST_SB_OUT_B16;
wire Tile_X05_Y0F_clk_out;
wire Tile_X05_Y0F_clk_pass_through_out_bot;
wire Tile_X05_Y0F_clk_pass_through_out_right;
wire [31:0] Tile_X05_Y0F_config_out_config_addr;
wire [31:0] Tile_X05_Y0F_config_out_config_data;
wire [0:0] Tile_X05_Y0F_config_out_read;
wire [0:0] Tile_X05_Y0F_config_out_write;
wire [8:0] Tile_X05_Y0F_hi_unq1;
wire [7:0] Tile_X05_Y0F_lo_unq1;
wire [31:0] Tile_X05_Y0F_read_config_data;
wire Tile_X05_Y0F_reset_out;
wire [0:0] Tile_X05_Y0F_stall_out;
wire [8:0] Tile_X05_Y0F_hi_out;
wire [7:0] Tile_X05_Y0F_lo_out;
wire [15:0] Tile_X05_Y0F_tile_id_in;
wire [0:0] Tile_X05_Y10_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y10_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y10_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y10_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y10_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y10_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y10_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y10_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y10_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y10_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y10_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y10_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y10_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y10_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y10_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y10_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y10_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y10_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y10_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y10_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y10_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y10_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y10_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y10_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y10_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y10_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y10_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y10_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y10_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y10_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y10_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y10_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X05_Y10_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X05_Y10_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X05_Y10_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y10_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y10_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X05_Y10_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X05_Y10_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X05_Y10_SB_T4_WEST_SB_OUT_B16;
wire Tile_X05_Y10_clk_out;
wire Tile_X05_Y10_clk_pass_through_out_bot;
wire Tile_X05_Y10_clk_pass_through_out_right;
wire [31:0] Tile_X05_Y10_config_out_config_addr;
wire [31:0] Tile_X05_Y10_config_out_config_data;
wire [0:0] Tile_X05_Y10_config_out_read;
wire [0:0] Tile_X05_Y10_config_out_write;
wire [8:0] Tile_X05_Y10_hi;
wire [7:0] Tile_X05_Y10_lo_unq1;
wire [31:0] Tile_X05_Y10_read_config_data;
wire Tile_X05_Y10_reset_out;
wire [0:0] Tile_X05_Y10_stall_out;
wire [7:0] Tile_X05_Y10_lo_out;
wire [15:0] Tile_X05_Y10_tile_id_in;
wire [0:0] Tile_X06_Y00_io2glb_1;
wire [0:0] Tile_X06_Y00_io2f_1;
wire [15:0] Tile_X06_Y00_io2glb_16;
wire [15:0] Tile_X06_Y00_io2f_16;
wire [8:0] Tile_X06_Y00_hi;
wire [7:0] Tile_X06_Y00_lo;
wire [0:0] Tile_X06_Y01_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y01_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y01_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y01_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y01_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y01_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y01_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y01_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y01_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y01_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y01_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y01_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y01_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y01_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y01_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y01_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y01_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y01_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y01_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y01_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y01_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y01_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y01_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y01_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y01_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y01_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y01_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y01_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y01_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y01_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y01_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y01_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y01_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y01_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y01_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y01_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y01_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y01_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y01_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y01_SB_T4_WEST_SB_OUT_B16;
wire Tile_X06_Y01_clk_out;
wire Tile_X06_Y01_clk_pass_through_out_bot;
wire Tile_X06_Y01_clk_pass_through_out_right;
wire [31:0] Tile_X06_Y01_config_out_config_addr;
wire [31:0] Tile_X06_Y01_config_out_config_data;
wire [0:0] Tile_X06_Y01_config_out_read;
wire [0:0] Tile_X06_Y01_config_out_write;
wire [8:0] Tile_X06_Y01_hi;
wire [7:0] Tile_X06_Y01_lo_unq1;
wire [31:0] Tile_X06_Y01_read_config_data;
wire Tile_X06_Y01_reset_out;
wire [0:0] Tile_X06_Y01_stall_out;
wire [7:0] Tile_X06_Y01_lo_out;
wire [15:0] Tile_X06_Y01_tile_id_in;
wire [0:0] Tile_X06_Y02_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y02_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y02_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y02_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y02_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y02_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y02_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y02_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y02_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y02_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y02_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y02_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y02_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y02_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y02_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y02_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y02_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y02_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y02_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y02_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y02_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y02_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y02_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y02_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y02_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y02_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y02_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y02_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y02_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y02_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y02_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y02_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y02_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y02_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y02_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y02_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y02_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y02_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y02_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y02_SB_T4_WEST_SB_OUT_B16;
wire Tile_X06_Y02_clk_out;
wire Tile_X06_Y02_clk_pass_through_out_bot;
wire Tile_X06_Y02_clk_pass_through_out_right;
wire [31:0] Tile_X06_Y02_config_out_config_addr;
wire [31:0] Tile_X06_Y02_config_out_config_data;
wire [0:0] Tile_X06_Y02_config_out_read;
wire [0:0] Tile_X06_Y02_config_out_write;
wire [8:0] Tile_X06_Y02_hi;
wire [7:0] Tile_X06_Y02_lo_unq1;
wire [31:0] Tile_X06_Y02_read_config_data;
wire Tile_X06_Y02_reset_out;
wire [0:0] Tile_X06_Y02_stall_out;
wire [7:0] Tile_X06_Y02_lo_out;
wire [15:0] Tile_X06_Y02_tile_id_in;
wire [0:0] Tile_X06_Y03_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y03_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y03_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y03_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y03_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y03_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y03_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y03_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y03_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y03_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y03_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y03_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y03_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y03_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y03_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y03_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y03_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y03_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y03_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y03_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y03_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y03_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y03_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y03_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y03_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y03_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y03_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y03_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y03_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y03_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y03_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y03_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y03_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y03_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y03_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y03_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y03_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y03_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y03_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y03_SB_T4_WEST_SB_OUT_B16;
wire Tile_X06_Y03_clk_out;
wire Tile_X06_Y03_clk_pass_through_out_bot;
wire Tile_X06_Y03_clk_pass_through_out_right;
wire [31:0] Tile_X06_Y03_config_out_config_addr;
wire [31:0] Tile_X06_Y03_config_out_config_data;
wire [0:0] Tile_X06_Y03_config_out_read;
wire [0:0] Tile_X06_Y03_config_out_write;
wire [8:0] Tile_X06_Y03_hi_unq1;
wire [7:0] Tile_X06_Y03_lo_unq1;
wire [31:0] Tile_X06_Y03_read_config_data;
wire Tile_X06_Y03_reset_out;
wire [0:0] Tile_X06_Y03_stall_out;
wire [8:0] Tile_X06_Y03_hi_out;
wire [7:0] Tile_X06_Y03_lo_out;
wire [15:0] Tile_X06_Y03_tile_id_in;
wire [0:0] Tile_X06_Y04_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y04_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y04_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y04_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y04_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y04_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y04_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y04_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y04_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y04_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y04_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y04_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y04_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y04_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y04_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y04_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y04_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y04_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y04_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y04_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y04_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y04_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y04_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y04_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y04_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y04_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y04_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y04_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y04_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y04_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y04_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y04_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y04_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y04_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y04_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y04_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y04_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y04_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y04_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y04_SB_T4_WEST_SB_OUT_B16;
wire Tile_X06_Y04_clk_out;
wire Tile_X06_Y04_clk_pass_through_out_bot;
wire Tile_X06_Y04_clk_pass_through_out_right;
wire [31:0] Tile_X06_Y04_config_out_config_addr;
wire [31:0] Tile_X06_Y04_config_out_config_data;
wire [0:0] Tile_X06_Y04_config_out_read;
wire [0:0] Tile_X06_Y04_config_out_write;
wire [8:0] Tile_X06_Y04_hi;
wire [7:0] Tile_X06_Y04_lo_unq1;
wire [31:0] Tile_X06_Y04_read_config_data;
wire Tile_X06_Y04_reset_out;
wire [0:0] Tile_X06_Y04_stall_out;
wire [7:0] Tile_X06_Y04_lo_out;
wire [15:0] Tile_X06_Y04_tile_id_in;
wire [0:0] Tile_X06_Y05_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y05_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y05_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y05_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y05_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y05_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y05_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y05_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y05_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y05_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y05_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y05_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y05_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y05_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y05_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y05_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y05_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y05_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y05_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y05_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y05_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y05_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y05_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y05_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y05_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y05_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y05_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y05_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y05_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y05_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y05_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y05_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y05_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y05_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y05_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y05_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y05_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y05_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y05_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y05_SB_T4_WEST_SB_OUT_B16;
wire Tile_X06_Y05_clk_out;
wire Tile_X06_Y05_clk_pass_through_out_bot;
wire Tile_X06_Y05_clk_pass_through_out_right;
wire [31:0] Tile_X06_Y05_config_out_config_addr;
wire [31:0] Tile_X06_Y05_config_out_config_data;
wire [0:0] Tile_X06_Y05_config_out_read;
wire [0:0] Tile_X06_Y05_config_out_write;
wire [8:0] Tile_X06_Y05_hi;
wire [7:0] Tile_X06_Y05_lo_unq1;
wire [31:0] Tile_X06_Y05_read_config_data;
wire Tile_X06_Y05_reset_out;
wire [0:0] Tile_X06_Y05_stall_out;
wire [7:0] Tile_X06_Y05_lo_out;
wire [15:0] Tile_X06_Y05_tile_id_in;
wire [0:0] Tile_X06_Y06_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y06_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y06_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y06_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y06_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y06_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y06_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y06_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y06_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y06_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y06_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y06_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y06_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y06_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y06_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y06_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y06_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y06_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y06_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y06_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y06_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y06_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y06_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y06_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y06_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y06_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y06_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y06_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y06_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y06_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y06_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y06_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y06_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y06_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y06_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y06_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y06_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y06_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y06_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y06_SB_T4_WEST_SB_OUT_B16;
wire Tile_X06_Y06_clk_out;
wire Tile_X06_Y06_clk_pass_through_out_bot;
wire Tile_X06_Y06_clk_pass_through_out_right;
wire [31:0] Tile_X06_Y06_config_out_config_addr;
wire [31:0] Tile_X06_Y06_config_out_config_data;
wire [0:0] Tile_X06_Y06_config_out_read;
wire [0:0] Tile_X06_Y06_config_out_write;
wire [8:0] Tile_X06_Y06_hi;
wire [7:0] Tile_X06_Y06_lo_unq1;
wire [31:0] Tile_X06_Y06_read_config_data;
wire Tile_X06_Y06_reset_out;
wire [0:0] Tile_X06_Y06_stall_out;
wire [7:0] Tile_X06_Y06_lo_out;
wire [15:0] Tile_X06_Y06_tile_id_in;
wire [0:0] Tile_X06_Y07_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y07_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y07_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y07_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y07_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y07_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y07_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y07_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y07_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y07_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y07_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y07_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y07_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y07_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y07_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y07_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y07_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y07_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y07_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y07_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y07_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y07_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y07_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y07_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y07_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y07_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y07_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y07_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y07_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y07_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y07_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y07_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y07_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y07_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y07_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y07_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y07_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y07_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y07_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y07_SB_T4_WEST_SB_OUT_B16;
wire Tile_X06_Y07_clk_out;
wire Tile_X06_Y07_clk_pass_through_out_bot;
wire Tile_X06_Y07_clk_pass_through_out_right;
wire [31:0] Tile_X06_Y07_config_out_config_addr;
wire [31:0] Tile_X06_Y07_config_out_config_data;
wire [0:0] Tile_X06_Y07_config_out_read;
wire [0:0] Tile_X06_Y07_config_out_write;
wire [8:0] Tile_X06_Y07_hi_unq1;
wire [7:0] Tile_X06_Y07_lo_unq1;
wire [31:0] Tile_X06_Y07_read_config_data;
wire Tile_X06_Y07_reset_out;
wire [0:0] Tile_X06_Y07_stall_out;
wire [8:0] Tile_X06_Y07_hi_out;
wire [7:0] Tile_X06_Y07_lo_out;
wire [15:0] Tile_X06_Y07_tile_id_in;
wire [0:0] Tile_X06_Y08_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y08_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y08_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y08_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y08_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y08_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y08_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y08_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y08_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y08_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y08_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y08_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y08_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y08_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y08_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y08_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y08_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y08_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y08_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y08_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y08_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y08_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y08_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y08_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y08_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y08_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y08_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y08_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y08_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y08_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y08_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y08_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y08_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y08_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y08_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y08_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y08_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y08_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y08_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y08_SB_T4_WEST_SB_OUT_B16;
wire Tile_X06_Y08_clk_out;
wire Tile_X06_Y08_clk_pass_through_out_bot;
wire Tile_X06_Y08_clk_pass_through_out_right;
wire [31:0] Tile_X06_Y08_config_out_config_addr;
wire [31:0] Tile_X06_Y08_config_out_config_data;
wire [0:0] Tile_X06_Y08_config_out_read;
wire [0:0] Tile_X06_Y08_config_out_write;
wire [8:0] Tile_X06_Y08_hi;
wire [7:0] Tile_X06_Y08_lo_unq1;
wire [31:0] Tile_X06_Y08_read_config_data;
wire Tile_X06_Y08_reset_out;
wire [0:0] Tile_X06_Y08_stall_out;
wire [7:0] Tile_X06_Y08_lo_out;
wire [15:0] Tile_X06_Y08_tile_id_in;
wire [0:0] Tile_X06_Y09_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y09_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y09_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y09_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y09_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y09_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y09_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y09_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y09_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y09_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y09_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y09_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y09_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y09_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y09_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y09_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y09_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y09_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y09_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y09_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y09_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y09_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y09_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y09_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y09_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y09_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y09_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y09_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y09_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y09_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y09_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y09_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y09_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y09_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y09_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y09_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y09_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y09_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y09_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y09_SB_T4_WEST_SB_OUT_B16;
wire Tile_X06_Y09_clk_out;
wire Tile_X06_Y09_clk_pass_through_out_bot;
wire Tile_X06_Y09_clk_pass_through_out_right;
wire [31:0] Tile_X06_Y09_config_out_config_addr;
wire [31:0] Tile_X06_Y09_config_out_config_data;
wire [0:0] Tile_X06_Y09_config_out_read;
wire [0:0] Tile_X06_Y09_config_out_write;
wire [8:0] Tile_X06_Y09_hi;
wire [7:0] Tile_X06_Y09_lo_unq1;
wire [31:0] Tile_X06_Y09_read_config_data;
wire Tile_X06_Y09_reset_out;
wire [0:0] Tile_X06_Y09_stall_out;
wire [7:0] Tile_X06_Y09_lo_out;
wire [15:0] Tile_X06_Y09_tile_id_in;
wire [0:0] Tile_X06_Y0A_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0A_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0A_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0A_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0A_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0A_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0A_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0A_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0A_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0A_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0A_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0A_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0A_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0A_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0A_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0A_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0A_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0A_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0A_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0A_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0A_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0A_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0A_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0A_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0A_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0A_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0A_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0A_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0A_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0A_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0A_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0A_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0A_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0A_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0A_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0A_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0A_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0A_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0A_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0A_SB_T4_WEST_SB_OUT_B16;
wire Tile_X06_Y0A_clk_out;
wire Tile_X06_Y0A_clk_pass_through_out_bot;
wire Tile_X06_Y0A_clk_pass_through_out_right;
wire [31:0] Tile_X06_Y0A_config_out_config_addr;
wire [31:0] Tile_X06_Y0A_config_out_config_data;
wire [0:0] Tile_X06_Y0A_config_out_read;
wire [0:0] Tile_X06_Y0A_config_out_write;
wire [8:0] Tile_X06_Y0A_hi;
wire [7:0] Tile_X06_Y0A_lo_unq1;
wire [31:0] Tile_X06_Y0A_read_config_data;
wire Tile_X06_Y0A_reset_out;
wire [0:0] Tile_X06_Y0A_stall_out;
wire [7:0] Tile_X06_Y0A_lo_out;
wire [15:0] Tile_X06_Y0A_tile_id_in;
wire [0:0] Tile_X06_Y0B_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0B_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0B_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0B_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0B_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0B_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0B_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0B_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0B_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0B_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0B_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0B_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0B_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0B_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0B_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0B_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0B_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0B_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0B_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0B_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0B_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0B_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0B_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0B_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0B_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0B_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0B_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0B_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0B_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0B_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0B_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0B_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0B_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0B_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0B_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0B_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0B_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0B_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0B_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0B_SB_T4_WEST_SB_OUT_B16;
wire Tile_X06_Y0B_clk_out;
wire Tile_X06_Y0B_clk_pass_through_out_bot;
wire Tile_X06_Y0B_clk_pass_through_out_right;
wire [31:0] Tile_X06_Y0B_config_out_config_addr;
wire [31:0] Tile_X06_Y0B_config_out_config_data;
wire [0:0] Tile_X06_Y0B_config_out_read;
wire [0:0] Tile_X06_Y0B_config_out_write;
wire [8:0] Tile_X06_Y0B_hi_unq1;
wire [7:0] Tile_X06_Y0B_lo_unq1;
wire [31:0] Tile_X06_Y0B_read_config_data;
wire Tile_X06_Y0B_reset_out;
wire [0:0] Tile_X06_Y0B_stall_out;
wire [8:0] Tile_X06_Y0B_hi_out;
wire [7:0] Tile_X06_Y0B_lo_out;
wire [15:0] Tile_X06_Y0B_tile_id_in;
wire [0:0] Tile_X06_Y0C_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0C_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0C_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0C_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0C_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0C_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0C_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0C_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0C_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0C_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0C_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0C_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0C_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0C_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0C_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0C_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0C_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0C_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0C_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0C_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0C_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0C_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0C_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0C_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0C_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0C_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0C_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0C_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0C_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0C_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0C_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0C_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0C_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0C_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0C_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0C_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0C_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0C_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0C_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0C_SB_T4_WEST_SB_OUT_B16;
wire Tile_X06_Y0C_clk_out;
wire Tile_X06_Y0C_clk_pass_through_out_bot;
wire Tile_X06_Y0C_clk_pass_through_out_right;
wire [31:0] Tile_X06_Y0C_config_out_config_addr;
wire [31:0] Tile_X06_Y0C_config_out_config_data;
wire [0:0] Tile_X06_Y0C_config_out_read;
wire [0:0] Tile_X06_Y0C_config_out_write;
wire [8:0] Tile_X06_Y0C_hi_unq1;
wire [7:0] Tile_X06_Y0C_lo_unq1;
wire [31:0] Tile_X06_Y0C_read_config_data;
wire Tile_X06_Y0C_reset_out;
wire [0:0] Tile_X06_Y0C_stall_out;
wire [8:0] Tile_X06_Y0C_hi_out;
wire [7:0] Tile_X06_Y0C_lo_out;
wire [15:0] Tile_X06_Y0C_tile_id_in;
wire [0:0] Tile_X06_Y0D_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0D_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0D_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0D_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0D_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0D_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0D_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0D_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0D_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0D_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0D_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0D_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0D_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0D_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0D_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0D_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0D_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0D_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0D_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0D_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0D_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0D_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0D_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0D_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0D_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0D_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0D_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0D_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0D_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0D_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0D_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0D_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0D_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0D_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0D_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0D_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0D_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0D_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0D_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0D_SB_T4_WEST_SB_OUT_B16;
wire Tile_X06_Y0D_clk_out;
wire Tile_X06_Y0D_clk_pass_through_out_bot;
wire Tile_X06_Y0D_clk_pass_through_out_right;
wire [31:0] Tile_X06_Y0D_config_out_config_addr;
wire [31:0] Tile_X06_Y0D_config_out_config_data;
wire [0:0] Tile_X06_Y0D_config_out_read;
wire [0:0] Tile_X06_Y0D_config_out_write;
wire [8:0] Tile_X06_Y0D_hi_unq1;
wire [7:0] Tile_X06_Y0D_lo_unq1;
wire [31:0] Tile_X06_Y0D_read_config_data;
wire Tile_X06_Y0D_reset_out;
wire [0:0] Tile_X06_Y0D_stall_out;
wire [8:0] Tile_X06_Y0D_hi_out;
wire [7:0] Tile_X06_Y0D_lo_out;
wire [15:0] Tile_X06_Y0D_tile_id_in;
wire [0:0] Tile_X06_Y0E_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0E_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0E_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0E_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0E_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0E_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0E_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0E_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0E_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0E_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0E_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0E_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0E_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0E_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0E_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0E_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0E_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0E_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0E_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0E_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0E_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0E_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0E_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0E_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0E_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0E_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0E_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0E_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0E_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0E_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0E_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0E_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0E_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0E_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0E_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0E_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0E_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0E_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0E_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0E_SB_T4_WEST_SB_OUT_B16;
wire Tile_X06_Y0E_clk_out;
wire Tile_X06_Y0E_clk_pass_through_out_bot;
wire Tile_X06_Y0E_clk_pass_through_out_right;
wire [31:0] Tile_X06_Y0E_config_out_config_addr;
wire [31:0] Tile_X06_Y0E_config_out_config_data;
wire [0:0] Tile_X06_Y0E_config_out_read;
wire [0:0] Tile_X06_Y0E_config_out_write;
wire [8:0] Tile_X06_Y0E_hi_unq1;
wire [7:0] Tile_X06_Y0E_lo_unq1;
wire [31:0] Tile_X06_Y0E_read_config_data;
wire Tile_X06_Y0E_reset_out;
wire [0:0] Tile_X06_Y0E_stall_out;
wire [8:0] Tile_X06_Y0E_hi_out;
wire [7:0] Tile_X06_Y0E_lo_out;
wire [15:0] Tile_X06_Y0E_tile_id_in;
wire [0:0] Tile_X06_Y0F_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0F_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0F_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0F_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0F_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0F_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0F_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0F_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0F_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0F_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0F_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0F_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0F_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0F_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0F_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0F_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0F_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0F_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0F_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0F_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0F_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0F_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0F_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0F_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0F_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0F_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0F_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0F_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0F_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0F_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0F_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0F_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0F_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0F_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y0F_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0F_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0F_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y0F_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y0F_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y0F_SB_T4_WEST_SB_OUT_B16;
wire Tile_X06_Y0F_clk_out;
wire Tile_X06_Y0F_clk_pass_through_out_bot;
wire Tile_X06_Y0F_clk_pass_through_out_right;
wire [31:0] Tile_X06_Y0F_config_out_config_addr;
wire [31:0] Tile_X06_Y0F_config_out_config_data;
wire [0:0] Tile_X06_Y0F_config_out_read;
wire [0:0] Tile_X06_Y0F_config_out_write;
wire [8:0] Tile_X06_Y0F_hi_unq1;
wire [7:0] Tile_X06_Y0F_lo_unq1;
wire [31:0] Tile_X06_Y0F_read_config_data;
wire Tile_X06_Y0F_reset_out;
wire [0:0] Tile_X06_Y0F_stall_out;
wire [8:0] Tile_X06_Y0F_hi_out;
wire [7:0] Tile_X06_Y0F_lo_out;
wire [15:0] Tile_X06_Y0F_tile_id_in;
wire [0:0] Tile_X06_Y10_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y10_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y10_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y10_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y10_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y10_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y10_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y10_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y10_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y10_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y10_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y10_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y10_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y10_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y10_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y10_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y10_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y10_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y10_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y10_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y10_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y10_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y10_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y10_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y10_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y10_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y10_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y10_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y10_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y10_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y10_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y10_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X06_Y10_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X06_Y10_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X06_Y10_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y10_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y10_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X06_Y10_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X06_Y10_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X06_Y10_SB_T4_WEST_SB_OUT_B16;
wire Tile_X06_Y10_clk_out;
wire Tile_X06_Y10_clk_pass_through_out_bot;
wire Tile_X06_Y10_clk_pass_through_out_right;
wire [31:0] Tile_X06_Y10_config_out_config_addr;
wire [31:0] Tile_X06_Y10_config_out_config_data;
wire [0:0] Tile_X06_Y10_config_out_read;
wire [0:0] Tile_X06_Y10_config_out_write;
wire [8:0] Tile_X06_Y10_hi;
wire [7:0] Tile_X06_Y10_lo_unq1;
wire [31:0] Tile_X06_Y10_read_config_data;
wire Tile_X06_Y10_reset_out;
wire [0:0] Tile_X06_Y10_stall_out;
wire [7:0] Tile_X06_Y10_lo_out;
wire [15:0] Tile_X06_Y10_tile_id_in;
wire [0:0] Tile_X07_Y00_io2glb_1;
wire [0:0] Tile_X07_Y00_io2f_1;
wire [15:0] Tile_X07_Y00_io2glb_16;
wire [15:0] Tile_X07_Y00_io2f_16;
wire [8:0] Tile_X07_Y00_hi;
wire [7:0] Tile_X07_Y00_lo;
wire [0:0] Tile_X07_Y01_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y01_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y01_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y01_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y01_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y01_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y01_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y01_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y01_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y01_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y01_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y01_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y01_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y01_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y01_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y01_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y01_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y01_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y01_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y01_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y01_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y01_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y01_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y01_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y01_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y01_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y01_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y01_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y01_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y01_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y01_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y01_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y01_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y01_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y01_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y01_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y01_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y01_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y01_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y01_SB_T4_WEST_SB_OUT_B16;
wire Tile_X07_Y01_clk_out;
wire [31:0] Tile_X07_Y01_config_out_config_addr;
wire [31:0] Tile_X07_Y01_config_out_config_data;
wire [0:0] Tile_X07_Y01_config_out_read;
wire [0:0] Tile_X07_Y01_config_out_write;
wire [8:0] Tile_X07_Y01_hi_unq1;
wire [7:0] Tile_X07_Y01_lo_unq1;
wire [31:0] Tile_X07_Y01_read_config_data;
wire Tile_X07_Y01_reset_out;
wire [0:0] Tile_X07_Y01_stall_out;
wire [8:0] Tile_X07_Y01_hi_out;
wire [7:0] Tile_X07_Y01_lo_out;
wire [15:0] Tile_X07_Y01_tile_id_in;
wire [0:0] Tile_X07_Y02_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y02_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y02_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y02_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y02_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y02_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y02_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y02_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y02_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y02_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y02_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y02_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y02_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y02_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y02_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y02_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y02_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y02_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y02_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y02_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y02_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y02_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y02_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y02_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y02_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y02_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y02_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y02_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y02_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y02_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y02_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y02_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y02_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y02_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y02_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y02_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y02_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y02_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y02_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y02_SB_T4_WEST_SB_OUT_B16;
wire Tile_X07_Y02_clk_out;
wire [31:0] Tile_X07_Y02_config_out_config_addr;
wire [31:0] Tile_X07_Y02_config_out_config_data;
wire [0:0] Tile_X07_Y02_config_out_read;
wire [0:0] Tile_X07_Y02_config_out_write;
wire [8:0] Tile_X07_Y02_hi_unq1;
wire [7:0] Tile_X07_Y02_lo_unq1;
wire [31:0] Tile_X07_Y02_read_config_data;
wire Tile_X07_Y02_reset_out;
wire [0:0] Tile_X07_Y02_stall_out;
wire [8:0] Tile_X07_Y02_hi_out;
wire [7:0] Tile_X07_Y02_lo_out;
wire [15:0] Tile_X07_Y02_tile_id_in;
wire [0:0] Tile_X07_Y03_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y03_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y03_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y03_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y03_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y03_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y03_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y03_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y03_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y03_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y03_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y03_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y03_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y03_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y03_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y03_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y03_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y03_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y03_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y03_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y03_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y03_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y03_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y03_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y03_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y03_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y03_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y03_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y03_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y03_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y03_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y03_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y03_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y03_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y03_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y03_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y03_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y03_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y03_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y03_SB_T4_WEST_SB_OUT_B16;
wire Tile_X07_Y03_clk_out;
wire [31:0] Tile_X07_Y03_config_out_config_addr;
wire [31:0] Tile_X07_Y03_config_out_config_data;
wire [0:0] Tile_X07_Y03_config_out_read;
wire [0:0] Tile_X07_Y03_config_out_write;
wire [8:0] Tile_X07_Y03_hi_unq1;
wire [7:0] Tile_X07_Y03_lo_unq1;
wire [31:0] Tile_X07_Y03_read_config_data;
wire Tile_X07_Y03_reset_out;
wire [0:0] Tile_X07_Y03_stall_out;
wire [8:0] Tile_X07_Y03_hi_out;
wire [7:0] Tile_X07_Y03_lo_out;
wire [15:0] Tile_X07_Y03_tile_id_in;
wire [0:0] Tile_X07_Y04_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y04_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y04_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y04_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y04_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y04_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y04_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y04_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y04_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y04_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y04_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y04_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y04_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y04_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y04_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y04_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y04_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y04_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y04_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y04_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y04_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y04_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y04_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y04_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y04_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y04_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y04_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y04_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y04_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y04_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y04_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y04_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y04_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y04_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y04_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y04_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y04_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y04_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y04_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y04_SB_T4_WEST_SB_OUT_B16;
wire Tile_X07_Y04_clk_out;
wire [31:0] Tile_X07_Y04_config_out_config_addr;
wire [31:0] Tile_X07_Y04_config_out_config_data;
wire [0:0] Tile_X07_Y04_config_out_read;
wire [0:0] Tile_X07_Y04_config_out_write;
wire [8:0] Tile_X07_Y04_hi_unq1;
wire [7:0] Tile_X07_Y04_lo_unq1;
wire [31:0] Tile_X07_Y04_read_config_data;
wire Tile_X07_Y04_reset_out;
wire [0:0] Tile_X07_Y04_stall_out;
wire [8:0] Tile_X07_Y04_hi_out;
wire [7:0] Tile_X07_Y04_lo_out;
wire [15:0] Tile_X07_Y04_tile_id_in;
wire [0:0] Tile_X07_Y05_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y05_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y05_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y05_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y05_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y05_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y05_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y05_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y05_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y05_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y05_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y05_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y05_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y05_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y05_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y05_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y05_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y05_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y05_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y05_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y05_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y05_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y05_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y05_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y05_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y05_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y05_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y05_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y05_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y05_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y05_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y05_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y05_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y05_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y05_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y05_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y05_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y05_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y05_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y05_SB_T4_WEST_SB_OUT_B16;
wire Tile_X07_Y05_clk_out;
wire [31:0] Tile_X07_Y05_config_out_config_addr;
wire [31:0] Tile_X07_Y05_config_out_config_data;
wire [0:0] Tile_X07_Y05_config_out_read;
wire [0:0] Tile_X07_Y05_config_out_write;
wire [8:0] Tile_X07_Y05_hi_unq1;
wire [7:0] Tile_X07_Y05_lo_unq1;
wire [31:0] Tile_X07_Y05_read_config_data;
wire Tile_X07_Y05_reset_out;
wire [0:0] Tile_X07_Y05_stall_out;
wire [8:0] Tile_X07_Y05_hi_out;
wire [7:0] Tile_X07_Y05_lo_out;
wire [15:0] Tile_X07_Y05_tile_id_in;
wire [0:0] Tile_X07_Y06_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y06_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y06_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y06_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y06_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y06_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y06_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y06_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y06_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y06_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y06_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y06_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y06_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y06_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y06_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y06_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y06_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y06_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y06_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y06_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y06_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y06_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y06_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y06_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y06_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y06_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y06_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y06_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y06_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y06_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y06_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y06_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y06_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y06_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y06_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y06_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y06_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y06_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y06_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y06_SB_T4_WEST_SB_OUT_B16;
wire Tile_X07_Y06_clk_out;
wire [31:0] Tile_X07_Y06_config_out_config_addr;
wire [31:0] Tile_X07_Y06_config_out_config_data;
wire [0:0] Tile_X07_Y06_config_out_read;
wire [0:0] Tile_X07_Y06_config_out_write;
wire [8:0] Tile_X07_Y06_hi_unq1;
wire [7:0] Tile_X07_Y06_lo_unq1;
wire [31:0] Tile_X07_Y06_read_config_data;
wire Tile_X07_Y06_reset_out;
wire [0:0] Tile_X07_Y06_stall_out;
wire [8:0] Tile_X07_Y06_hi_out;
wire [7:0] Tile_X07_Y06_lo_out;
wire [15:0] Tile_X07_Y06_tile_id_in;
wire [0:0] Tile_X07_Y07_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y07_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y07_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y07_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y07_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y07_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y07_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y07_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y07_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y07_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y07_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y07_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y07_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y07_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y07_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y07_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y07_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y07_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y07_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y07_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y07_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y07_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y07_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y07_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y07_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y07_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y07_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y07_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y07_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y07_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y07_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y07_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y07_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y07_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y07_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y07_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y07_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y07_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y07_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y07_SB_T4_WEST_SB_OUT_B16;
wire Tile_X07_Y07_clk_out;
wire [31:0] Tile_X07_Y07_config_out_config_addr;
wire [31:0] Tile_X07_Y07_config_out_config_data;
wire [0:0] Tile_X07_Y07_config_out_read;
wire [0:0] Tile_X07_Y07_config_out_write;
wire [8:0] Tile_X07_Y07_hi_unq1;
wire [7:0] Tile_X07_Y07_lo_unq1;
wire [31:0] Tile_X07_Y07_read_config_data;
wire Tile_X07_Y07_reset_out;
wire [0:0] Tile_X07_Y07_stall_out;
wire [8:0] Tile_X07_Y07_hi_out;
wire [7:0] Tile_X07_Y07_lo_out;
wire [15:0] Tile_X07_Y07_tile_id_in;
wire [0:0] Tile_X07_Y08_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y08_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y08_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y08_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y08_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y08_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y08_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y08_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y08_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y08_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y08_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y08_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y08_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y08_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y08_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y08_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y08_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y08_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y08_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y08_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y08_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y08_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y08_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y08_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y08_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y08_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y08_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y08_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y08_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y08_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y08_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y08_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y08_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y08_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y08_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y08_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y08_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y08_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y08_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y08_SB_T4_WEST_SB_OUT_B16;
wire Tile_X07_Y08_clk_out;
wire [31:0] Tile_X07_Y08_config_out_config_addr;
wire [31:0] Tile_X07_Y08_config_out_config_data;
wire [0:0] Tile_X07_Y08_config_out_read;
wire [0:0] Tile_X07_Y08_config_out_write;
wire [8:0] Tile_X07_Y08_hi_unq1;
wire [7:0] Tile_X07_Y08_lo_unq1;
wire [31:0] Tile_X07_Y08_read_config_data;
wire Tile_X07_Y08_reset_out;
wire [0:0] Tile_X07_Y08_stall_out;
wire [8:0] Tile_X07_Y08_hi_out;
wire [7:0] Tile_X07_Y08_lo_out;
wire [15:0] Tile_X07_Y08_tile_id_in;
wire [0:0] Tile_X07_Y09_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y09_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y09_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y09_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y09_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y09_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y09_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y09_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y09_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y09_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y09_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y09_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y09_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y09_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y09_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y09_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y09_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y09_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y09_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y09_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y09_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y09_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y09_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y09_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y09_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y09_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y09_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y09_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y09_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y09_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y09_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y09_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y09_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y09_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y09_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y09_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y09_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y09_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y09_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y09_SB_T4_WEST_SB_OUT_B16;
wire Tile_X07_Y09_clk_out;
wire [31:0] Tile_X07_Y09_config_out_config_addr;
wire [31:0] Tile_X07_Y09_config_out_config_data;
wire [0:0] Tile_X07_Y09_config_out_read;
wire [0:0] Tile_X07_Y09_config_out_write;
wire [8:0] Tile_X07_Y09_hi_unq1;
wire [7:0] Tile_X07_Y09_lo_unq1;
wire [31:0] Tile_X07_Y09_read_config_data;
wire Tile_X07_Y09_reset_out;
wire [0:0] Tile_X07_Y09_stall_out;
wire [8:0] Tile_X07_Y09_hi_out;
wire [7:0] Tile_X07_Y09_lo_out;
wire [15:0] Tile_X07_Y09_tile_id_in;
wire [0:0] Tile_X07_Y0A_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0A_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0A_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0A_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0A_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0A_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0A_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0A_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0A_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0A_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0A_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0A_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0A_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0A_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0A_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0A_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0A_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0A_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0A_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0A_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0A_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0A_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0A_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0A_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0A_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0A_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0A_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0A_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0A_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0A_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0A_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0A_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0A_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0A_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0A_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0A_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0A_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0A_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0A_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0A_SB_T4_WEST_SB_OUT_B16;
wire Tile_X07_Y0A_clk_out;
wire [31:0] Tile_X07_Y0A_config_out_config_addr;
wire [31:0] Tile_X07_Y0A_config_out_config_data;
wire [0:0] Tile_X07_Y0A_config_out_read;
wire [0:0] Tile_X07_Y0A_config_out_write;
wire [8:0] Tile_X07_Y0A_hi_unq1;
wire [7:0] Tile_X07_Y0A_lo_unq1;
wire [31:0] Tile_X07_Y0A_read_config_data;
wire Tile_X07_Y0A_reset_out;
wire [0:0] Tile_X07_Y0A_stall_out;
wire [8:0] Tile_X07_Y0A_hi_out;
wire [7:0] Tile_X07_Y0A_lo_out;
wire [15:0] Tile_X07_Y0A_tile_id_in;
wire [0:0] Tile_X07_Y0B_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0B_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0B_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0B_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0B_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0B_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0B_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0B_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0B_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0B_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0B_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0B_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0B_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0B_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0B_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0B_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0B_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0B_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0B_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0B_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0B_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0B_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0B_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0B_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0B_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0B_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0B_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0B_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0B_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0B_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0B_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0B_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0B_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0B_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0B_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0B_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0B_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0B_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0B_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0B_SB_T4_WEST_SB_OUT_B16;
wire Tile_X07_Y0B_clk_out;
wire [31:0] Tile_X07_Y0B_config_out_config_addr;
wire [31:0] Tile_X07_Y0B_config_out_config_data;
wire [0:0] Tile_X07_Y0B_config_out_read;
wire [0:0] Tile_X07_Y0B_config_out_write;
wire [8:0] Tile_X07_Y0B_hi_unq1;
wire [7:0] Tile_X07_Y0B_lo_unq1;
wire [31:0] Tile_X07_Y0B_read_config_data;
wire Tile_X07_Y0B_reset_out;
wire [0:0] Tile_X07_Y0B_stall_out;
wire [8:0] Tile_X07_Y0B_hi_out;
wire [7:0] Tile_X07_Y0B_lo_out;
wire [15:0] Tile_X07_Y0B_tile_id_in;
wire [0:0] Tile_X07_Y0C_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0C_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0C_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0C_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0C_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0C_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0C_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0C_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0C_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0C_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0C_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0C_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0C_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0C_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0C_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0C_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0C_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0C_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0C_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0C_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0C_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0C_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0C_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0C_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0C_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0C_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0C_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0C_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0C_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0C_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0C_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0C_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0C_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0C_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0C_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0C_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0C_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0C_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0C_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0C_SB_T4_WEST_SB_OUT_B16;
wire Tile_X07_Y0C_clk_out;
wire [31:0] Tile_X07_Y0C_config_out_config_addr;
wire [31:0] Tile_X07_Y0C_config_out_config_data;
wire [0:0] Tile_X07_Y0C_config_out_read;
wire [0:0] Tile_X07_Y0C_config_out_write;
wire [8:0] Tile_X07_Y0C_hi_unq1;
wire [7:0] Tile_X07_Y0C_lo_unq1;
wire [31:0] Tile_X07_Y0C_read_config_data;
wire Tile_X07_Y0C_reset_out;
wire [0:0] Tile_X07_Y0C_stall_out;
wire [8:0] Tile_X07_Y0C_hi_out;
wire [7:0] Tile_X07_Y0C_lo_out;
wire [15:0] Tile_X07_Y0C_tile_id_in;
wire [0:0] Tile_X07_Y0D_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0D_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0D_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0D_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0D_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0D_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0D_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0D_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0D_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0D_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0D_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0D_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0D_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0D_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0D_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0D_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0D_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0D_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0D_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0D_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0D_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0D_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0D_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0D_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0D_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0D_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0D_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0D_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0D_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0D_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0D_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0D_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0D_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0D_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0D_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0D_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0D_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0D_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0D_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0D_SB_T4_WEST_SB_OUT_B16;
wire Tile_X07_Y0D_clk_out;
wire [31:0] Tile_X07_Y0D_config_out_config_addr;
wire [31:0] Tile_X07_Y0D_config_out_config_data;
wire [0:0] Tile_X07_Y0D_config_out_read;
wire [0:0] Tile_X07_Y0D_config_out_write;
wire [8:0] Tile_X07_Y0D_hi_unq1;
wire [7:0] Tile_X07_Y0D_lo_unq1;
wire [31:0] Tile_X07_Y0D_read_config_data;
wire Tile_X07_Y0D_reset_out;
wire [0:0] Tile_X07_Y0D_stall_out;
wire [8:0] Tile_X07_Y0D_hi_out;
wire [7:0] Tile_X07_Y0D_lo_out;
wire [15:0] Tile_X07_Y0D_tile_id_in;
wire [0:0] Tile_X07_Y0E_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0E_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0E_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0E_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0E_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0E_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0E_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0E_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0E_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0E_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0E_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0E_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0E_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0E_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0E_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0E_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0E_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0E_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0E_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0E_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0E_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0E_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0E_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0E_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0E_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0E_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0E_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0E_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0E_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0E_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0E_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0E_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0E_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0E_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0E_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0E_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0E_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0E_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0E_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0E_SB_T4_WEST_SB_OUT_B16;
wire Tile_X07_Y0E_clk_out;
wire [31:0] Tile_X07_Y0E_config_out_config_addr;
wire [31:0] Tile_X07_Y0E_config_out_config_data;
wire [0:0] Tile_X07_Y0E_config_out_read;
wire [0:0] Tile_X07_Y0E_config_out_write;
wire [8:0] Tile_X07_Y0E_hi_unq1;
wire [7:0] Tile_X07_Y0E_lo_unq1;
wire [31:0] Tile_X07_Y0E_read_config_data;
wire Tile_X07_Y0E_reset_out;
wire [0:0] Tile_X07_Y0E_stall_out;
wire [8:0] Tile_X07_Y0E_hi_out;
wire [7:0] Tile_X07_Y0E_lo_out;
wire [15:0] Tile_X07_Y0E_tile_id_in;
wire [0:0] Tile_X07_Y0F_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0F_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0F_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0F_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0F_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0F_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0F_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0F_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0F_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0F_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0F_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0F_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0F_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0F_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0F_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0F_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0F_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0F_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0F_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0F_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0F_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0F_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0F_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0F_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0F_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0F_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0F_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0F_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0F_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0F_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0F_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0F_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0F_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0F_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y0F_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0F_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0F_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y0F_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y0F_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y0F_SB_T4_WEST_SB_OUT_B16;
wire Tile_X07_Y0F_clk_out;
wire [31:0] Tile_X07_Y0F_config_out_config_addr;
wire [31:0] Tile_X07_Y0F_config_out_config_data;
wire [0:0] Tile_X07_Y0F_config_out_read;
wire [0:0] Tile_X07_Y0F_config_out_write;
wire [8:0] Tile_X07_Y0F_hi_unq1;
wire [7:0] Tile_X07_Y0F_lo_unq1;
wire [31:0] Tile_X07_Y0F_read_config_data;
wire Tile_X07_Y0F_reset_out;
wire [0:0] Tile_X07_Y0F_stall_out;
wire [8:0] Tile_X07_Y0F_hi_out;
wire [7:0] Tile_X07_Y0F_lo_out;
wire [15:0] Tile_X07_Y0F_tile_id_in;
wire [0:0] Tile_X07_Y10_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y10_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y10_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y10_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y10_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y10_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y10_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y10_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y10_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y10_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y10_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y10_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y10_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y10_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y10_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y10_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y10_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y10_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y10_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y10_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y10_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y10_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y10_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y10_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y10_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y10_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y10_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y10_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y10_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y10_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y10_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y10_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X07_Y10_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X07_Y10_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X07_Y10_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y10_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y10_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X07_Y10_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X07_Y10_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X07_Y10_SB_T4_WEST_SB_OUT_B16;
wire Tile_X07_Y10_clk_out;
wire [31:0] Tile_X07_Y10_config_out_config_addr;
wire [31:0] Tile_X07_Y10_config_out_config_data;
wire [0:0] Tile_X07_Y10_config_out_read;
wire [0:0] Tile_X07_Y10_config_out_write;
wire [8:0] Tile_X07_Y10_hi_unq1;
wire [7:0] Tile_X07_Y10_lo_unq1;
wire [31:0] Tile_X07_Y10_read_config_data;
wire Tile_X07_Y10_reset_out;
wire [0:0] Tile_X07_Y10_stall_out;
wire [8:0] Tile_X07_Y10_hi_out;
wire [7:0] Tile_X07_Y10_lo_out;
wire [15:0] Tile_X07_Y10_tile_id_in;
wire [0:0] Tile_X08_Y00_io2glb_1;
wire [0:0] Tile_X08_Y00_io2f_1;
wire [15:0] Tile_X08_Y00_io2glb_16;
wire [15:0] Tile_X08_Y00_io2f_16;
wire [8:0] Tile_X08_Y00_hi;
wire [7:0] Tile_X08_Y00_lo;
wire [0:0] Tile_X08_Y01_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y01_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y01_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y01_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y01_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y01_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y01_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y01_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y01_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y01_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y01_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y01_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y01_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y01_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y01_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y01_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y01_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y01_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y01_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y01_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y01_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y01_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y01_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y01_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y01_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y01_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y01_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y01_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y01_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y01_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y01_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y01_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y01_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y01_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y01_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y01_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y01_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y01_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y01_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y01_SB_T4_WEST_SB_OUT_B16;
wire Tile_X08_Y01_clk_out;
wire Tile_X08_Y01_clk_pass_through_out_bot;
wire Tile_X08_Y01_clk_pass_through_out_right;
wire [31:0] Tile_X08_Y01_config_out_config_addr;
wire [31:0] Tile_X08_Y01_config_out_config_data;
wire [0:0] Tile_X08_Y01_config_out_read;
wire [0:0] Tile_X08_Y01_config_out_write;
wire [8:0] Tile_X08_Y01_hi;
wire [7:0] Tile_X08_Y01_lo_unq1;
wire [31:0] Tile_X08_Y01_read_config_data;
wire Tile_X08_Y01_reset_out;
wire [0:0] Tile_X08_Y01_stall_out;
wire [7:0] Tile_X08_Y01_lo_out;
wire [15:0] Tile_X08_Y01_tile_id_in;
wire [0:0] Tile_X08_Y02_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y02_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y02_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y02_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y02_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y02_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y02_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y02_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y02_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y02_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y02_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y02_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y02_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y02_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y02_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y02_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y02_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y02_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y02_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y02_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y02_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y02_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y02_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y02_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y02_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y02_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y02_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y02_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y02_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y02_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y02_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y02_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y02_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y02_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y02_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y02_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y02_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y02_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y02_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y02_SB_T4_WEST_SB_OUT_B16;
wire Tile_X08_Y02_clk_out;
wire Tile_X08_Y02_clk_pass_through_out_bot;
wire Tile_X08_Y02_clk_pass_through_out_right;
wire [31:0] Tile_X08_Y02_config_out_config_addr;
wire [31:0] Tile_X08_Y02_config_out_config_data;
wire [0:0] Tile_X08_Y02_config_out_read;
wire [0:0] Tile_X08_Y02_config_out_write;
wire [8:0] Tile_X08_Y02_hi;
wire [7:0] Tile_X08_Y02_lo_unq1;
wire [31:0] Tile_X08_Y02_read_config_data;
wire Tile_X08_Y02_reset_out;
wire [0:0] Tile_X08_Y02_stall_out;
wire [7:0] Tile_X08_Y02_lo_out;
wire [15:0] Tile_X08_Y02_tile_id_in;
wire [0:0] Tile_X08_Y03_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y03_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y03_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y03_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y03_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y03_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y03_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y03_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y03_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y03_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y03_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y03_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y03_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y03_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y03_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y03_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y03_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y03_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y03_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y03_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y03_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y03_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y03_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y03_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y03_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y03_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y03_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y03_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y03_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y03_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y03_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y03_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y03_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y03_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y03_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y03_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y03_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y03_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y03_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y03_SB_T4_WEST_SB_OUT_B16;
wire Tile_X08_Y03_clk_out;
wire Tile_X08_Y03_clk_pass_through_out_bot;
wire Tile_X08_Y03_clk_pass_through_out_right;
wire [31:0] Tile_X08_Y03_config_out_config_addr;
wire [31:0] Tile_X08_Y03_config_out_config_data;
wire [0:0] Tile_X08_Y03_config_out_read;
wire [0:0] Tile_X08_Y03_config_out_write;
wire [8:0] Tile_X08_Y03_hi_unq1;
wire [7:0] Tile_X08_Y03_lo_unq1;
wire [31:0] Tile_X08_Y03_read_config_data;
wire Tile_X08_Y03_reset_out;
wire [0:0] Tile_X08_Y03_stall_out;
wire [8:0] Tile_X08_Y03_hi_out;
wire [7:0] Tile_X08_Y03_lo_out;
wire [15:0] Tile_X08_Y03_tile_id_in;
wire [0:0] Tile_X08_Y04_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y04_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y04_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y04_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y04_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y04_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y04_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y04_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y04_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y04_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y04_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y04_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y04_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y04_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y04_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y04_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y04_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y04_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y04_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y04_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y04_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y04_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y04_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y04_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y04_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y04_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y04_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y04_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y04_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y04_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y04_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y04_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y04_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y04_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y04_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y04_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y04_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y04_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y04_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y04_SB_T4_WEST_SB_OUT_B16;
wire Tile_X08_Y04_clk_out;
wire Tile_X08_Y04_clk_pass_through_out_bot;
wire Tile_X08_Y04_clk_pass_through_out_right;
wire [31:0] Tile_X08_Y04_config_out_config_addr;
wire [31:0] Tile_X08_Y04_config_out_config_data;
wire [0:0] Tile_X08_Y04_config_out_read;
wire [0:0] Tile_X08_Y04_config_out_write;
wire [8:0] Tile_X08_Y04_hi;
wire [7:0] Tile_X08_Y04_lo_unq1;
wire [31:0] Tile_X08_Y04_read_config_data;
wire Tile_X08_Y04_reset_out;
wire [0:0] Tile_X08_Y04_stall_out;
wire [7:0] Tile_X08_Y04_lo_out;
wire [15:0] Tile_X08_Y04_tile_id_in;
wire [0:0] Tile_X08_Y05_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y05_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y05_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y05_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y05_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y05_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y05_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y05_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y05_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y05_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y05_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y05_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y05_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y05_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y05_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y05_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y05_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y05_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y05_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y05_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y05_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y05_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y05_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y05_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y05_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y05_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y05_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y05_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y05_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y05_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y05_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y05_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y05_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y05_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y05_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y05_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y05_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y05_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y05_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y05_SB_T4_WEST_SB_OUT_B16;
wire Tile_X08_Y05_clk_out;
wire Tile_X08_Y05_clk_pass_through_out_bot;
wire Tile_X08_Y05_clk_pass_through_out_right;
wire [31:0] Tile_X08_Y05_config_out_config_addr;
wire [31:0] Tile_X08_Y05_config_out_config_data;
wire [0:0] Tile_X08_Y05_config_out_read;
wire [0:0] Tile_X08_Y05_config_out_write;
wire [8:0] Tile_X08_Y05_hi;
wire [7:0] Tile_X08_Y05_lo_unq1;
wire [31:0] Tile_X08_Y05_read_config_data;
wire Tile_X08_Y05_reset_out;
wire [0:0] Tile_X08_Y05_stall_out;
wire [7:0] Tile_X08_Y05_lo_out;
wire [15:0] Tile_X08_Y05_tile_id_in;
wire [0:0] Tile_X08_Y06_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y06_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y06_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y06_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y06_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y06_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y06_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y06_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y06_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y06_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y06_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y06_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y06_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y06_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y06_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y06_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y06_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y06_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y06_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y06_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y06_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y06_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y06_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y06_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y06_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y06_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y06_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y06_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y06_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y06_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y06_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y06_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y06_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y06_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y06_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y06_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y06_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y06_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y06_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y06_SB_T4_WEST_SB_OUT_B16;
wire Tile_X08_Y06_clk_out;
wire Tile_X08_Y06_clk_pass_through_out_bot;
wire Tile_X08_Y06_clk_pass_through_out_right;
wire [31:0] Tile_X08_Y06_config_out_config_addr;
wire [31:0] Tile_X08_Y06_config_out_config_data;
wire [0:0] Tile_X08_Y06_config_out_read;
wire [0:0] Tile_X08_Y06_config_out_write;
wire [8:0] Tile_X08_Y06_hi;
wire [7:0] Tile_X08_Y06_lo_unq1;
wire [31:0] Tile_X08_Y06_read_config_data;
wire Tile_X08_Y06_reset_out;
wire [0:0] Tile_X08_Y06_stall_out;
wire [7:0] Tile_X08_Y06_lo_out;
wire [15:0] Tile_X08_Y06_tile_id_in;
wire [0:0] Tile_X08_Y07_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y07_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y07_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y07_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y07_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y07_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y07_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y07_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y07_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y07_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y07_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y07_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y07_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y07_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y07_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y07_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y07_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y07_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y07_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y07_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y07_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y07_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y07_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y07_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y07_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y07_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y07_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y07_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y07_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y07_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y07_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y07_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y07_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y07_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y07_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y07_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y07_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y07_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y07_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y07_SB_T4_WEST_SB_OUT_B16;
wire Tile_X08_Y07_clk_out;
wire Tile_X08_Y07_clk_pass_through_out_bot;
wire Tile_X08_Y07_clk_pass_through_out_right;
wire [31:0] Tile_X08_Y07_config_out_config_addr;
wire [31:0] Tile_X08_Y07_config_out_config_data;
wire [0:0] Tile_X08_Y07_config_out_read;
wire [0:0] Tile_X08_Y07_config_out_write;
wire [8:0] Tile_X08_Y07_hi_unq1;
wire [7:0] Tile_X08_Y07_lo_unq1;
wire [31:0] Tile_X08_Y07_read_config_data;
wire Tile_X08_Y07_reset_out;
wire [0:0] Tile_X08_Y07_stall_out;
wire [8:0] Tile_X08_Y07_hi_out;
wire [7:0] Tile_X08_Y07_lo_out;
wire [15:0] Tile_X08_Y07_tile_id_in;
wire [0:0] Tile_X08_Y08_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y08_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y08_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y08_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y08_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y08_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y08_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y08_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y08_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y08_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y08_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y08_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y08_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y08_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y08_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y08_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y08_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y08_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y08_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y08_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y08_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y08_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y08_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y08_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y08_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y08_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y08_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y08_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y08_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y08_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y08_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y08_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y08_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y08_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y08_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y08_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y08_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y08_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y08_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y08_SB_T4_WEST_SB_OUT_B16;
wire Tile_X08_Y08_clk_out;
wire Tile_X08_Y08_clk_pass_through_out_bot;
wire Tile_X08_Y08_clk_pass_through_out_right;
wire [31:0] Tile_X08_Y08_config_out_config_addr;
wire [31:0] Tile_X08_Y08_config_out_config_data;
wire [0:0] Tile_X08_Y08_config_out_read;
wire [0:0] Tile_X08_Y08_config_out_write;
wire [8:0] Tile_X08_Y08_hi;
wire [7:0] Tile_X08_Y08_lo_unq1;
wire [31:0] Tile_X08_Y08_read_config_data;
wire Tile_X08_Y08_reset_out;
wire [0:0] Tile_X08_Y08_stall_out;
wire [7:0] Tile_X08_Y08_lo_out;
wire [15:0] Tile_X08_Y08_tile_id_in;
wire [0:0] Tile_X08_Y09_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y09_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y09_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y09_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y09_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y09_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y09_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y09_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y09_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y09_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y09_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y09_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y09_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y09_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y09_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y09_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y09_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y09_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y09_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y09_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y09_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y09_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y09_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y09_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y09_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y09_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y09_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y09_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y09_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y09_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y09_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y09_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y09_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y09_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y09_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y09_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y09_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y09_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y09_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y09_SB_T4_WEST_SB_OUT_B16;
wire Tile_X08_Y09_clk_out;
wire Tile_X08_Y09_clk_pass_through_out_bot;
wire Tile_X08_Y09_clk_pass_through_out_right;
wire [31:0] Tile_X08_Y09_config_out_config_addr;
wire [31:0] Tile_X08_Y09_config_out_config_data;
wire [0:0] Tile_X08_Y09_config_out_read;
wire [0:0] Tile_X08_Y09_config_out_write;
wire [8:0] Tile_X08_Y09_hi;
wire [7:0] Tile_X08_Y09_lo_unq1;
wire [31:0] Tile_X08_Y09_read_config_data;
wire Tile_X08_Y09_reset_out;
wire [0:0] Tile_X08_Y09_stall_out;
wire [7:0] Tile_X08_Y09_lo_out;
wire [15:0] Tile_X08_Y09_tile_id_in;
wire [0:0] Tile_X08_Y0A_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0A_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0A_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0A_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0A_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0A_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0A_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0A_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0A_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0A_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0A_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0A_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0A_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0A_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0A_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0A_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0A_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0A_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0A_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0A_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0A_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0A_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0A_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0A_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0A_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0A_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0A_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0A_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0A_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0A_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0A_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0A_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0A_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0A_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0A_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0A_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0A_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0A_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0A_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0A_SB_T4_WEST_SB_OUT_B16;
wire Tile_X08_Y0A_clk_out;
wire Tile_X08_Y0A_clk_pass_through_out_bot;
wire Tile_X08_Y0A_clk_pass_through_out_right;
wire [31:0] Tile_X08_Y0A_config_out_config_addr;
wire [31:0] Tile_X08_Y0A_config_out_config_data;
wire [0:0] Tile_X08_Y0A_config_out_read;
wire [0:0] Tile_X08_Y0A_config_out_write;
wire [8:0] Tile_X08_Y0A_hi;
wire [7:0] Tile_X08_Y0A_lo_unq1;
wire [31:0] Tile_X08_Y0A_read_config_data;
wire Tile_X08_Y0A_reset_out;
wire [0:0] Tile_X08_Y0A_stall_out;
wire [7:0] Tile_X08_Y0A_lo_out;
wire [15:0] Tile_X08_Y0A_tile_id_in;
wire [0:0] Tile_X08_Y0B_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0B_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0B_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0B_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0B_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0B_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0B_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0B_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0B_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0B_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0B_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0B_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0B_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0B_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0B_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0B_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0B_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0B_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0B_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0B_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0B_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0B_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0B_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0B_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0B_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0B_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0B_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0B_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0B_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0B_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0B_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0B_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0B_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0B_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0B_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0B_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0B_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0B_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0B_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0B_SB_T4_WEST_SB_OUT_B16;
wire Tile_X08_Y0B_clk_out;
wire Tile_X08_Y0B_clk_pass_through_out_bot;
wire Tile_X08_Y0B_clk_pass_through_out_right;
wire [31:0] Tile_X08_Y0B_config_out_config_addr;
wire [31:0] Tile_X08_Y0B_config_out_config_data;
wire [0:0] Tile_X08_Y0B_config_out_read;
wire [0:0] Tile_X08_Y0B_config_out_write;
wire [8:0] Tile_X08_Y0B_hi_unq1;
wire [7:0] Tile_X08_Y0B_lo_unq1;
wire [31:0] Tile_X08_Y0B_read_config_data;
wire Tile_X08_Y0B_reset_out;
wire [0:0] Tile_X08_Y0B_stall_out;
wire [8:0] Tile_X08_Y0B_hi_out;
wire [7:0] Tile_X08_Y0B_lo_out;
wire [15:0] Tile_X08_Y0B_tile_id_in;
wire [0:0] Tile_X08_Y0C_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0C_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0C_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0C_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0C_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0C_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0C_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0C_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0C_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0C_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0C_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0C_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0C_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0C_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0C_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0C_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0C_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0C_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0C_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0C_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0C_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0C_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0C_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0C_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0C_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0C_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0C_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0C_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0C_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0C_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0C_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0C_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0C_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0C_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0C_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0C_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0C_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0C_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0C_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0C_SB_T4_WEST_SB_OUT_B16;
wire Tile_X08_Y0C_clk_out;
wire Tile_X08_Y0C_clk_pass_through_out_bot;
wire Tile_X08_Y0C_clk_pass_through_out_right;
wire [31:0] Tile_X08_Y0C_config_out_config_addr;
wire [31:0] Tile_X08_Y0C_config_out_config_data;
wire [0:0] Tile_X08_Y0C_config_out_read;
wire [0:0] Tile_X08_Y0C_config_out_write;
wire [8:0] Tile_X08_Y0C_hi_unq1;
wire [7:0] Tile_X08_Y0C_lo_unq1;
wire [31:0] Tile_X08_Y0C_read_config_data;
wire Tile_X08_Y0C_reset_out;
wire [0:0] Tile_X08_Y0C_stall_out;
wire [8:0] Tile_X08_Y0C_hi_out;
wire [7:0] Tile_X08_Y0C_lo_out;
wire [15:0] Tile_X08_Y0C_tile_id_in;
wire [0:0] Tile_X08_Y0D_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0D_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0D_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0D_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0D_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0D_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0D_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0D_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0D_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0D_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0D_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0D_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0D_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0D_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0D_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0D_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0D_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0D_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0D_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0D_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0D_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0D_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0D_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0D_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0D_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0D_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0D_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0D_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0D_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0D_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0D_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0D_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0D_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0D_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0D_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0D_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0D_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0D_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0D_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0D_SB_T4_WEST_SB_OUT_B16;
wire Tile_X08_Y0D_clk_out;
wire Tile_X08_Y0D_clk_pass_through_out_bot;
wire Tile_X08_Y0D_clk_pass_through_out_right;
wire [31:0] Tile_X08_Y0D_config_out_config_addr;
wire [31:0] Tile_X08_Y0D_config_out_config_data;
wire [0:0] Tile_X08_Y0D_config_out_read;
wire [0:0] Tile_X08_Y0D_config_out_write;
wire [8:0] Tile_X08_Y0D_hi_unq1;
wire [7:0] Tile_X08_Y0D_lo_unq1;
wire [31:0] Tile_X08_Y0D_read_config_data;
wire Tile_X08_Y0D_reset_out;
wire [0:0] Tile_X08_Y0D_stall_out;
wire [8:0] Tile_X08_Y0D_hi_out;
wire [7:0] Tile_X08_Y0D_lo_out;
wire [15:0] Tile_X08_Y0D_tile_id_in;
wire [0:0] Tile_X08_Y0E_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0E_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0E_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0E_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0E_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0E_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0E_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0E_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0E_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0E_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0E_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0E_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0E_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0E_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0E_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0E_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0E_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0E_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0E_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0E_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0E_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0E_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0E_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0E_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0E_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0E_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0E_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0E_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0E_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0E_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0E_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0E_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0E_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0E_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0E_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0E_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0E_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0E_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0E_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0E_SB_T4_WEST_SB_OUT_B16;
wire Tile_X08_Y0E_clk_out;
wire Tile_X08_Y0E_clk_pass_through_out_bot;
wire Tile_X08_Y0E_clk_pass_through_out_right;
wire [31:0] Tile_X08_Y0E_config_out_config_addr;
wire [31:0] Tile_X08_Y0E_config_out_config_data;
wire [0:0] Tile_X08_Y0E_config_out_read;
wire [0:0] Tile_X08_Y0E_config_out_write;
wire [8:0] Tile_X08_Y0E_hi_unq1;
wire [7:0] Tile_X08_Y0E_lo_unq1;
wire [31:0] Tile_X08_Y0E_read_config_data;
wire Tile_X08_Y0E_reset_out;
wire [0:0] Tile_X08_Y0E_stall_out;
wire [8:0] Tile_X08_Y0E_hi_out;
wire [7:0] Tile_X08_Y0E_lo_out;
wire [15:0] Tile_X08_Y0E_tile_id_in;
wire [0:0] Tile_X08_Y0F_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0F_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0F_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0F_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0F_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0F_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0F_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0F_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0F_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0F_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0F_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0F_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0F_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0F_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0F_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0F_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0F_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0F_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0F_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0F_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0F_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0F_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0F_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0F_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0F_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0F_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0F_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0F_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0F_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0F_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0F_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0F_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0F_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0F_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y0F_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0F_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0F_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y0F_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y0F_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y0F_SB_T4_WEST_SB_OUT_B16;
wire Tile_X08_Y0F_clk_out;
wire Tile_X08_Y0F_clk_pass_through_out_bot;
wire Tile_X08_Y0F_clk_pass_through_out_right;
wire [31:0] Tile_X08_Y0F_config_out_config_addr;
wire [31:0] Tile_X08_Y0F_config_out_config_data;
wire [0:0] Tile_X08_Y0F_config_out_read;
wire [0:0] Tile_X08_Y0F_config_out_write;
wire [8:0] Tile_X08_Y0F_hi_unq1;
wire [7:0] Tile_X08_Y0F_lo_unq1;
wire [31:0] Tile_X08_Y0F_read_config_data;
wire Tile_X08_Y0F_reset_out;
wire [0:0] Tile_X08_Y0F_stall_out;
wire [8:0] Tile_X08_Y0F_hi_out;
wire [7:0] Tile_X08_Y0F_lo_out;
wire [15:0] Tile_X08_Y0F_tile_id_in;
wire [0:0] Tile_X08_Y10_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y10_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y10_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y10_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y10_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y10_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y10_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y10_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y10_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y10_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y10_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y10_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y10_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y10_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y10_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y10_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y10_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y10_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y10_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y10_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y10_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y10_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y10_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y10_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y10_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y10_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y10_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y10_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y10_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y10_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y10_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y10_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X08_Y10_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X08_Y10_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X08_Y10_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y10_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y10_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X08_Y10_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X08_Y10_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X08_Y10_SB_T4_WEST_SB_OUT_B16;
wire Tile_X08_Y10_clk_out;
wire Tile_X08_Y10_clk_pass_through_out_bot;
wire Tile_X08_Y10_clk_pass_through_out_right;
wire [31:0] Tile_X08_Y10_config_out_config_addr;
wire [31:0] Tile_X08_Y10_config_out_config_data;
wire [0:0] Tile_X08_Y10_config_out_read;
wire [0:0] Tile_X08_Y10_config_out_write;
wire [8:0] Tile_X08_Y10_hi;
wire [7:0] Tile_X08_Y10_lo_unq1;
wire [31:0] Tile_X08_Y10_read_config_data;
wire Tile_X08_Y10_reset_out;
wire [0:0] Tile_X08_Y10_stall_out;
wire [7:0] Tile_X08_Y10_lo_out;
wire [15:0] Tile_X08_Y10_tile_id_in;
wire [0:0] Tile_X09_Y00_io2glb_1;
wire [0:0] Tile_X09_Y00_io2f_1;
wire [15:0] Tile_X09_Y00_io2glb_16;
wire [15:0] Tile_X09_Y00_io2f_16;
wire [8:0] Tile_X09_Y00_hi;
wire [7:0] Tile_X09_Y00_lo;
wire [0:0] Tile_X09_Y01_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y01_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y01_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y01_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y01_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y01_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y01_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y01_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y01_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y01_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y01_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y01_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y01_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y01_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y01_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y01_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y01_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y01_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y01_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y01_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y01_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y01_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y01_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y01_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y01_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y01_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y01_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y01_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y01_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y01_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y01_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y01_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y01_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y01_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y01_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y01_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y01_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y01_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y01_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y01_SB_T4_WEST_SB_OUT_B16;
wire Tile_X09_Y01_clk_out;
wire Tile_X09_Y01_clk_pass_through_out_bot;
wire Tile_X09_Y01_clk_pass_through_out_right;
wire [31:0] Tile_X09_Y01_config_out_config_addr;
wire [31:0] Tile_X09_Y01_config_out_config_data;
wire [0:0] Tile_X09_Y01_config_out_read;
wire [0:0] Tile_X09_Y01_config_out_write;
wire [8:0] Tile_X09_Y01_hi;
wire [7:0] Tile_X09_Y01_lo_unq1;
wire [31:0] Tile_X09_Y01_read_config_data;
wire Tile_X09_Y01_reset_out;
wire [0:0] Tile_X09_Y01_stall_out;
wire [7:0] Tile_X09_Y01_lo_out;
wire [15:0] Tile_X09_Y01_tile_id_in;
wire [0:0] Tile_X09_Y02_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y02_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y02_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y02_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y02_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y02_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y02_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y02_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y02_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y02_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y02_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y02_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y02_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y02_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y02_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y02_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y02_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y02_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y02_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y02_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y02_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y02_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y02_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y02_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y02_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y02_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y02_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y02_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y02_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y02_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y02_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y02_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y02_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y02_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y02_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y02_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y02_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y02_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y02_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y02_SB_T4_WEST_SB_OUT_B16;
wire Tile_X09_Y02_clk_out;
wire Tile_X09_Y02_clk_pass_through_out_bot;
wire Tile_X09_Y02_clk_pass_through_out_right;
wire [31:0] Tile_X09_Y02_config_out_config_addr;
wire [31:0] Tile_X09_Y02_config_out_config_data;
wire [0:0] Tile_X09_Y02_config_out_read;
wire [0:0] Tile_X09_Y02_config_out_write;
wire [8:0] Tile_X09_Y02_hi;
wire [7:0] Tile_X09_Y02_lo_unq1;
wire [31:0] Tile_X09_Y02_read_config_data;
wire Tile_X09_Y02_reset_out;
wire [0:0] Tile_X09_Y02_stall_out;
wire [7:0] Tile_X09_Y02_lo_out;
wire [15:0] Tile_X09_Y02_tile_id_in;
wire [0:0] Tile_X09_Y03_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y03_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y03_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y03_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y03_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y03_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y03_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y03_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y03_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y03_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y03_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y03_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y03_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y03_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y03_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y03_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y03_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y03_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y03_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y03_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y03_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y03_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y03_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y03_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y03_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y03_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y03_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y03_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y03_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y03_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y03_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y03_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y03_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y03_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y03_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y03_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y03_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y03_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y03_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y03_SB_T4_WEST_SB_OUT_B16;
wire Tile_X09_Y03_clk_out;
wire Tile_X09_Y03_clk_pass_through_out_bot;
wire Tile_X09_Y03_clk_pass_through_out_right;
wire [31:0] Tile_X09_Y03_config_out_config_addr;
wire [31:0] Tile_X09_Y03_config_out_config_data;
wire [0:0] Tile_X09_Y03_config_out_read;
wire [0:0] Tile_X09_Y03_config_out_write;
wire [8:0] Tile_X09_Y03_hi_unq1;
wire [7:0] Tile_X09_Y03_lo_unq1;
wire [31:0] Tile_X09_Y03_read_config_data;
wire Tile_X09_Y03_reset_out;
wire [0:0] Tile_X09_Y03_stall_out;
wire [8:0] Tile_X09_Y03_hi_out;
wire [7:0] Tile_X09_Y03_lo_out;
wire [15:0] Tile_X09_Y03_tile_id_in;
wire [0:0] Tile_X09_Y04_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y04_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y04_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y04_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y04_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y04_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y04_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y04_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y04_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y04_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y04_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y04_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y04_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y04_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y04_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y04_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y04_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y04_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y04_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y04_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y04_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y04_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y04_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y04_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y04_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y04_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y04_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y04_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y04_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y04_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y04_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y04_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y04_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y04_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y04_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y04_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y04_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y04_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y04_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y04_SB_T4_WEST_SB_OUT_B16;
wire Tile_X09_Y04_clk_out;
wire Tile_X09_Y04_clk_pass_through_out_bot;
wire Tile_X09_Y04_clk_pass_through_out_right;
wire [31:0] Tile_X09_Y04_config_out_config_addr;
wire [31:0] Tile_X09_Y04_config_out_config_data;
wire [0:0] Tile_X09_Y04_config_out_read;
wire [0:0] Tile_X09_Y04_config_out_write;
wire [8:0] Tile_X09_Y04_hi;
wire [7:0] Tile_X09_Y04_lo_unq1;
wire [31:0] Tile_X09_Y04_read_config_data;
wire Tile_X09_Y04_reset_out;
wire [0:0] Tile_X09_Y04_stall_out;
wire [7:0] Tile_X09_Y04_lo_out;
wire [15:0] Tile_X09_Y04_tile_id_in;
wire [0:0] Tile_X09_Y05_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y05_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y05_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y05_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y05_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y05_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y05_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y05_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y05_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y05_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y05_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y05_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y05_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y05_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y05_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y05_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y05_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y05_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y05_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y05_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y05_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y05_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y05_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y05_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y05_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y05_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y05_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y05_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y05_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y05_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y05_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y05_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y05_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y05_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y05_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y05_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y05_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y05_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y05_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y05_SB_T4_WEST_SB_OUT_B16;
wire Tile_X09_Y05_clk_out;
wire Tile_X09_Y05_clk_pass_through_out_bot;
wire Tile_X09_Y05_clk_pass_through_out_right;
wire [31:0] Tile_X09_Y05_config_out_config_addr;
wire [31:0] Tile_X09_Y05_config_out_config_data;
wire [0:0] Tile_X09_Y05_config_out_read;
wire [0:0] Tile_X09_Y05_config_out_write;
wire [8:0] Tile_X09_Y05_hi;
wire [7:0] Tile_X09_Y05_lo_unq1;
wire [31:0] Tile_X09_Y05_read_config_data;
wire Tile_X09_Y05_reset_out;
wire [0:0] Tile_X09_Y05_stall_out;
wire [7:0] Tile_X09_Y05_lo_out;
wire [15:0] Tile_X09_Y05_tile_id_in;
wire [0:0] Tile_X09_Y06_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y06_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y06_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y06_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y06_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y06_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y06_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y06_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y06_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y06_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y06_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y06_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y06_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y06_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y06_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y06_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y06_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y06_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y06_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y06_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y06_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y06_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y06_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y06_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y06_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y06_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y06_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y06_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y06_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y06_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y06_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y06_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y06_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y06_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y06_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y06_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y06_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y06_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y06_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y06_SB_T4_WEST_SB_OUT_B16;
wire Tile_X09_Y06_clk_out;
wire Tile_X09_Y06_clk_pass_through_out_bot;
wire Tile_X09_Y06_clk_pass_through_out_right;
wire [31:0] Tile_X09_Y06_config_out_config_addr;
wire [31:0] Tile_X09_Y06_config_out_config_data;
wire [0:0] Tile_X09_Y06_config_out_read;
wire [0:0] Tile_X09_Y06_config_out_write;
wire [8:0] Tile_X09_Y06_hi;
wire [7:0] Tile_X09_Y06_lo_unq1;
wire [31:0] Tile_X09_Y06_read_config_data;
wire Tile_X09_Y06_reset_out;
wire [0:0] Tile_X09_Y06_stall_out;
wire [7:0] Tile_X09_Y06_lo_out;
wire [15:0] Tile_X09_Y06_tile_id_in;
wire [0:0] Tile_X09_Y07_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y07_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y07_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y07_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y07_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y07_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y07_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y07_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y07_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y07_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y07_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y07_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y07_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y07_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y07_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y07_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y07_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y07_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y07_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y07_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y07_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y07_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y07_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y07_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y07_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y07_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y07_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y07_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y07_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y07_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y07_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y07_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y07_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y07_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y07_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y07_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y07_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y07_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y07_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y07_SB_T4_WEST_SB_OUT_B16;
wire Tile_X09_Y07_clk_out;
wire Tile_X09_Y07_clk_pass_through_out_bot;
wire Tile_X09_Y07_clk_pass_through_out_right;
wire [31:0] Tile_X09_Y07_config_out_config_addr;
wire [31:0] Tile_X09_Y07_config_out_config_data;
wire [0:0] Tile_X09_Y07_config_out_read;
wire [0:0] Tile_X09_Y07_config_out_write;
wire [8:0] Tile_X09_Y07_hi_unq1;
wire [7:0] Tile_X09_Y07_lo_unq1;
wire [31:0] Tile_X09_Y07_read_config_data;
wire Tile_X09_Y07_reset_out;
wire [0:0] Tile_X09_Y07_stall_out;
wire [8:0] Tile_X09_Y07_hi_out;
wire [7:0] Tile_X09_Y07_lo_out;
wire [15:0] Tile_X09_Y07_tile_id_in;
wire [0:0] Tile_X09_Y08_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y08_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y08_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y08_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y08_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y08_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y08_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y08_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y08_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y08_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y08_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y08_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y08_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y08_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y08_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y08_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y08_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y08_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y08_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y08_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y08_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y08_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y08_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y08_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y08_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y08_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y08_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y08_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y08_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y08_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y08_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y08_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y08_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y08_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y08_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y08_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y08_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y08_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y08_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y08_SB_T4_WEST_SB_OUT_B16;
wire Tile_X09_Y08_clk_out;
wire Tile_X09_Y08_clk_pass_through_out_bot;
wire Tile_X09_Y08_clk_pass_through_out_right;
wire [31:0] Tile_X09_Y08_config_out_config_addr;
wire [31:0] Tile_X09_Y08_config_out_config_data;
wire [0:0] Tile_X09_Y08_config_out_read;
wire [0:0] Tile_X09_Y08_config_out_write;
wire [8:0] Tile_X09_Y08_hi;
wire [7:0] Tile_X09_Y08_lo_unq1;
wire [31:0] Tile_X09_Y08_read_config_data;
wire Tile_X09_Y08_reset_out;
wire [0:0] Tile_X09_Y08_stall_out;
wire [7:0] Tile_X09_Y08_lo_out;
wire [15:0] Tile_X09_Y08_tile_id_in;
wire [0:0] Tile_X09_Y09_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y09_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y09_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y09_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y09_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y09_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y09_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y09_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y09_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y09_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y09_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y09_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y09_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y09_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y09_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y09_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y09_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y09_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y09_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y09_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y09_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y09_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y09_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y09_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y09_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y09_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y09_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y09_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y09_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y09_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y09_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y09_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y09_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y09_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y09_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y09_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y09_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y09_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y09_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y09_SB_T4_WEST_SB_OUT_B16;
wire Tile_X09_Y09_clk_out;
wire Tile_X09_Y09_clk_pass_through_out_bot;
wire Tile_X09_Y09_clk_pass_through_out_right;
wire [31:0] Tile_X09_Y09_config_out_config_addr;
wire [31:0] Tile_X09_Y09_config_out_config_data;
wire [0:0] Tile_X09_Y09_config_out_read;
wire [0:0] Tile_X09_Y09_config_out_write;
wire [8:0] Tile_X09_Y09_hi;
wire [7:0] Tile_X09_Y09_lo_unq1;
wire [31:0] Tile_X09_Y09_read_config_data;
wire Tile_X09_Y09_reset_out;
wire [0:0] Tile_X09_Y09_stall_out;
wire [7:0] Tile_X09_Y09_lo_out;
wire [15:0] Tile_X09_Y09_tile_id_in;
wire [0:0] Tile_X09_Y0A_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0A_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0A_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0A_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0A_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0A_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0A_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0A_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0A_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0A_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0A_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0A_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0A_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0A_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0A_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0A_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0A_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0A_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0A_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0A_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0A_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0A_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0A_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0A_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0A_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0A_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0A_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0A_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0A_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0A_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0A_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0A_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0A_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0A_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0A_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0A_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0A_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0A_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0A_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0A_SB_T4_WEST_SB_OUT_B16;
wire Tile_X09_Y0A_clk_out;
wire Tile_X09_Y0A_clk_pass_through_out_bot;
wire Tile_X09_Y0A_clk_pass_through_out_right;
wire [31:0] Tile_X09_Y0A_config_out_config_addr;
wire [31:0] Tile_X09_Y0A_config_out_config_data;
wire [0:0] Tile_X09_Y0A_config_out_read;
wire [0:0] Tile_X09_Y0A_config_out_write;
wire [8:0] Tile_X09_Y0A_hi;
wire [7:0] Tile_X09_Y0A_lo_unq1;
wire [31:0] Tile_X09_Y0A_read_config_data;
wire Tile_X09_Y0A_reset_out;
wire [0:0] Tile_X09_Y0A_stall_out;
wire [7:0] Tile_X09_Y0A_lo_out;
wire [15:0] Tile_X09_Y0A_tile_id_in;
wire [0:0] Tile_X09_Y0B_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0B_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0B_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0B_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0B_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0B_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0B_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0B_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0B_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0B_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0B_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0B_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0B_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0B_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0B_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0B_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0B_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0B_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0B_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0B_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0B_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0B_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0B_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0B_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0B_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0B_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0B_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0B_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0B_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0B_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0B_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0B_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0B_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0B_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0B_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0B_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0B_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0B_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0B_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0B_SB_T4_WEST_SB_OUT_B16;
wire Tile_X09_Y0B_clk_out;
wire Tile_X09_Y0B_clk_pass_through_out_bot;
wire Tile_X09_Y0B_clk_pass_through_out_right;
wire [31:0] Tile_X09_Y0B_config_out_config_addr;
wire [31:0] Tile_X09_Y0B_config_out_config_data;
wire [0:0] Tile_X09_Y0B_config_out_read;
wire [0:0] Tile_X09_Y0B_config_out_write;
wire [8:0] Tile_X09_Y0B_hi_unq1;
wire [7:0] Tile_X09_Y0B_lo_unq1;
wire [31:0] Tile_X09_Y0B_read_config_data;
wire Tile_X09_Y0B_reset_out;
wire [0:0] Tile_X09_Y0B_stall_out;
wire [8:0] Tile_X09_Y0B_hi_out;
wire [7:0] Tile_X09_Y0B_lo_out;
wire [15:0] Tile_X09_Y0B_tile_id_in;
wire [0:0] Tile_X09_Y0C_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0C_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0C_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0C_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0C_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0C_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0C_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0C_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0C_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0C_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0C_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0C_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0C_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0C_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0C_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0C_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0C_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0C_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0C_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0C_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0C_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0C_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0C_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0C_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0C_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0C_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0C_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0C_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0C_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0C_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0C_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0C_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0C_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0C_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0C_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0C_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0C_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0C_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0C_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0C_SB_T4_WEST_SB_OUT_B16;
wire Tile_X09_Y0C_clk_out;
wire Tile_X09_Y0C_clk_pass_through_out_bot;
wire Tile_X09_Y0C_clk_pass_through_out_right;
wire [31:0] Tile_X09_Y0C_config_out_config_addr;
wire [31:0] Tile_X09_Y0C_config_out_config_data;
wire [0:0] Tile_X09_Y0C_config_out_read;
wire [0:0] Tile_X09_Y0C_config_out_write;
wire [8:0] Tile_X09_Y0C_hi_unq1;
wire [7:0] Tile_X09_Y0C_lo_unq1;
wire [31:0] Tile_X09_Y0C_read_config_data;
wire Tile_X09_Y0C_reset_out;
wire [0:0] Tile_X09_Y0C_stall_out;
wire [8:0] Tile_X09_Y0C_hi_out;
wire [7:0] Tile_X09_Y0C_lo_out;
wire [15:0] Tile_X09_Y0C_tile_id_in;
wire [0:0] Tile_X09_Y0D_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0D_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0D_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0D_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0D_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0D_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0D_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0D_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0D_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0D_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0D_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0D_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0D_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0D_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0D_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0D_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0D_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0D_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0D_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0D_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0D_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0D_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0D_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0D_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0D_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0D_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0D_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0D_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0D_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0D_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0D_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0D_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0D_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0D_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0D_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0D_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0D_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0D_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0D_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0D_SB_T4_WEST_SB_OUT_B16;
wire Tile_X09_Y0D_clk_out;
wire Tile_X09_Y0D_clk_pass_through_out_bot;
wire Tile_X09_Y0D_clk_pass_through_out_right;
wire [31:0] Tile_X09_Y0D_config_out_config_addr;
wire [31:0] Tile_X09_Y0D_config_out_config_data;
wire [0:0] Tile_X09_Y0D_config_out_read;
wire [0:0] Tile_X09_Y0D_config_out_write;
wire [8:0] Tile_X09_Y0D_hi_unq1;
wire [7:0] Tile_X09_Y0D_lo_unq1;
wire [31:0] Tile_X09_Y0D_read_config_data;
wire Tile_X09_Y0D_reset_out;
wire [0:0] Tile_X09_Y0D_stall_out;
wire [8:0] Tile_X09_Y0D_hi_out;
wire [7:0] Tile_X09_Y0D_lo_out;
wire [15:0] Tile_X09_Y0D_tile_id_in;
wire [0:0] Tile_X09_Y0E_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0E_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0E_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0E_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0E_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0E_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0E_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0E_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0E_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0E_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0E_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0E_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0E_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0E_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0E_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0E_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0E_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0E_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0E_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0E_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0E_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0E_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0E_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0E_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0E_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0E_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0E_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0E_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0E_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0E_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0E_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0E_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0E_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0E_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0E_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0E_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0E_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0E_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0E_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0E_SB_T4_WEST_SB_OUT_B16;
wire Tile_X09_Y0E_clk_out;
wire Tile_X09_Y0E_clk_pass_through_out_bot;
wire Tile_X09_Y0E_clk_pass_through_out_right;
wire [31:0] Tile_X09_Y0E_config_out_config_addr;
wire [31:0] Tile_X09_Y0E_config_out_config_data;
wire [0:0] Tile_X09_Y0E_config_out_read;
wire [0:0] Tile_X09_Y0E_config_out_write;
wire [8:0] Tile_X09_Y0E_hi_unq1;
wire [7:0] Tile_X09_Y0E_lo_unq1;
wire [31:0] Tile_X09_Y0E_read_config_data;
wire Tile_X09_Y0E_reset_out;
wire [0:0] Tile_X09_Y0E_stall_out;
wire [8:0] Tile_X09_Y0E_hi_out;
wire [7:0] Tile_X09_Y0E_lo_out;
wire [15:0] Tile_X09_Y0E_tile_id_in;
wire [0:0] Tile_X09_Y0F_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0F_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0F_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0F_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0F_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0F_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0F_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0F_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0F_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0F_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0F_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0F_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0F_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0F_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0F_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0F_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0F_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0F_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0F_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0F_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0F_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0F_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0F_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0F_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0F_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0F_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0F_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0F_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0F_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0F_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0F_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0F_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0F_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0F_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y0F_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0F_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0F_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y0F_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y0F_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y0F_SB_T4_WEST_SB_OUT_B16;
wire Tile_X09_Y0F_clk_out;
wire Tile_X09_Y0F_clk_pass_through_out_bot;
wire Tile_X09_Y0F_clk_pass_through_out_right;
wire [31:0] Tile_X09_Y0F_config_out_config_addr;
wire [31:0] Tile_X09_Y0F_config_out_config_data;
wire [0:0] Tile_X09_Y0F_config_out_read;
wire [0:0] Tile_X09_Y0F_config_out_write;
wire [8:0] Tile_X09_Y0F_hi_unq1;
wire [7:0] Tile_X09_Y0F_lo_unq1;
wire [31:0] Tile_X09_Y0F_read_config_data;
wire Tile_X09_Y0F_reset_out;
wire [0:0] Tile_X09_Y0F_stall_out;
wire [8:0] Tile_X09_Y0F_hi_out;
wire [7:0] Tile_X09_Y0F_lo_out;
wire [15:0] Tile_X09_Y0F_tile_id_in;
wire [0:0] Tile_X09_Y10_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y10_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y10_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y10_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y10_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y10_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y10_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y10_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y10_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y10_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y10_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y10_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y10_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y10_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y10_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y10_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y10_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y10_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y10_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y10_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y10_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y10_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y10_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y10_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y10_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y10_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y10_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y10_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y10_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y10_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y10_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y10_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X09_Y10_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X09_Y10_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X09_Y10_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y10_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y10_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X09_Y10_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X09_Y10_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X09_Y10_SB_T4_WEST_SB_OUT_B16;
wire Tile_X09_Y10_clk_out;
wire Tile_X09_Y10_clk_pass_through_out_bot;
wire Tile_X09_Y10_clk_pass_through_out_right;
wire [31:0] Tile_X09_Y10_config_out_config_addr;
wire [31:0] Tile_X09_Y10_config_out_config_data;
wire [0:0] Tile_X09_Y10_config_out_read;
wire [0:0] Tile_X09_Y10_config_out_write;
wire [8:0] Tile_X09_Y10_hi;
wire [7:0] Tile_X09_Y10_lo_unq1;
wire [31:0] Tile_X09_Y10_read_config_data;
wire Tile_X09_Y10_reset_out;
wire [0:0] Tile_X09_Y10_stall_out;
wire [7:0] Tile_X09_Y10_lo_out;
wire [15:0] Tile_X09_Y10_tile_id_in;
wire [0:0] Tile_X0A_Y00_io2glb_1;
wire [0:0] Tile_X0A_Y00_io2f_1;
wire [15:0] Tile_X0A_Y00_io2glb_16;
wire [15:0] Tile_X0A_Y00_io2f_16;
wire [8:0] Tile_X0A_Y00_hi;
wire [7:0] Tile_X0A_Y00_lo;
wire [0:0] Tile_X0A_Y01_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y01_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y01_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y01_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y01_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y01_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y01_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y01_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y01_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y01_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y01_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y01_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y01_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y01_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y01_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y01_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y01_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y01_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y01_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y01_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y01_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y01_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y01_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y01_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y01_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y01_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y01_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y01_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y01_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y01_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y01_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y01_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y01_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y01_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y01_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y01_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y01_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y01_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y01_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y01_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0A_Y01_clk_out;
wire Tile_X0A_Y01_clk_pass_through_out_bot;
wire Tile_X0A_Y01_clk_pass_through_out_right;
wire [31:0] Tile_X0A_Y01_config_out_config_addr;
wire [31:0] Tile_X0A_Y01_config_out_config_data;
wire [0:0] Tile_X0A_Y01_config_out_read;
wire [0:0] Tile_X0A_Y01_config_out_write;
wire [8:0] Tile_X0A_Y01_hi;
wire [7:0] Tile_X0A_Y01_lo_unq1;
wire [31:0] Tile_X0A_Y01_read_config_data;
wire Tile_X0A_Y01_reset_out;
wire [0:0] Tile_X0A_Y01_stall_out;
wire [7:0] Tile_X0A_Y01_lo_out;
wire [15:0] Tile_X0A_Y01_tile_id_in;
wire [0:0] Tile_X0A_Y02_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y02_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y02_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y02_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y02_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y02_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y02_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y02_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y02_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y02_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y02_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y02_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y02_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y02_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y02_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y02_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y02_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y02_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y02_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y02_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y02_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y02_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y02_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y02_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y02_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y02_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y02_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y02_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y02_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y02_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y02_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y02_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y02_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y02_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y02_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y02_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y02_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y02_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y02_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y02_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0A_Y02_clk_out;
wire Tile_X0A_Y02_clk_pass_through_out_bot;
wire Tile_X0A_Y02_clk_pass_through_out_right;
wire [31:0] Tile_X0A_Y02_config_out_config_addr;
wire [31:0] Tile_X0A_Y02_config_out_config_data;
wire [0:0] Tile_X0A_Y02_config_out_read;
wire [0:0] Tile_X0A_Y02_config_out_write;
wire [8:0] Tile_X0A_Y02_hi;
wire [7:0] Tile_X0A_Y02_lo_unq1;
wire [31:0] Tile_X0A_Y02_read_config_data;
wire Tile_X0A_Y02_reset_out;
wire [0:0] Tile_X0A_Y02_stall_out;
wire [7:0] Tile_X0A_Y02_lo_out;
wire [15:0] Tile_X0A_Y02_tile_id_in;
wire [0:0] Tile_X0A_Y03_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y03_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y03_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y03_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y03_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y03_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y03_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y03_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y03_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y03_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y03_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y03_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y03_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y03_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y03_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y03_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y03_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y03_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y03_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y03_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y03_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y03_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y03_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y03_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y03_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y03_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y03_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y03_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y03_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y03_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y03_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y03_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y03_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y03_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y03_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y03_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y03_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y03_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y03_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y03_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0A_Y03_clk_out;
wire Tile_X0A_Y03_clk_pass_through_out_bot;
wire Tile_X0A_Y03_clk_pass_through_out_right;
wire [31:0] Tile_X0A_Y03_config_out_config_addr;
wire [31:0] Tile_X0A_Y03_config_out_config_data;
wire [0:0] Tile_X0A_Y03_config_out_read;
wire [0:0] Tile_X0A_Y03_config_out_write;
wire [8:0] Tile_X0A_Y03_hi_unq1;
wire [7:0] Tile_X0A_Y03_lo_unq1;
wire [31:0] Tile_X0A_Y03_read_config_data;
wire Tile_X0A_Y03_reset_out;
wire [0:0] Tile_X0A_Y03_stall_out;
wire [8:0] Tile_X0A_Y03_hi_out;
wire [7:0] Tile_X0A_Y03_lo_out;
wire [15:0] Tile_X0A_Y03_tile_id_in;
wire [0:0] Tile_X0A_Y04_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y04_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y04_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y04_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y04_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y04_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y04_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y04_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y04_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y04_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y04_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y04_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y04_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y04_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y04_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y04_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y04_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y04_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y04_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y04_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y04_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y04_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y04_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y04_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y04_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y04_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y04_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y04_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y04_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y04_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y04_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y04_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y04_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y04_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y04_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y04_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y04_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y04_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y04_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y04_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0A_Y04_clk_out;
wire Tile_X0A_Y04_clk_pass_through_out_bot;
wire Tile_X0A_Y04_clk_pass_through_out_right;
wire [31:0] Tile_X0A_Y04_config_out_config_addr;
wire [31:0] Tile_X0A_Y04_config_out_config_data;
wire [0:0] Tile_X0A_Y04_config_out_read;
wire [0:0] Tile_X0A_Y04_config_out_write;
wire [8:0] Tile_X0A_Y04_hi;
wire [7:0] Tile_X0A_Y04_lo_unq1;
wire [31:0] Tile_X0A_Y04_read_config_data;
wire Tile_X0A_Y04_reset_out;
wire [0:0] Tile_X0A_Y04_stall_out;
wire [7:0] Tile_X0A_Y04_lo_out;
wire [15:0] Tile_X0A_Y04_tile_id_in;
wire [0:0] Tile_X0A_Y05_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y05_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y05_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y05_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y05_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y05_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y05_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y05_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y05_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y05_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y05_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y05_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y05_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y05_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y05_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y05_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y05_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y05_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y05_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y05_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y05_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y05_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y05_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y05_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y05_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y05_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y05_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y05_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y05_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y05_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y05_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y05_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y05_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y05_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y05_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y05_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y05_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y05_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y05_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y05_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0A_Y05_clk_out;
wire Tile_X0A_Y05_clk_pass_through_out_bot;
wire Tile_X0A_Y05_clk_pass_through_out_right;
wire [31:0] Tile_X0A_Y05_config_out_config_addr;
wire [31:0] Tile_X0A_Y05_config_out_config_data;
wire [0:0] Tile_X0A_Y05_config_out_read;
wire [0:0] Tile_X0A_Y05_config_out_write;
wire [8:0] Tile_X0A_Y05_hi;
wire [7:0] Tile_X0A_Y05_lo_unq1;
wire [31:0] Tile_X0A_Y05_read_config_data;
wire Tile_X0A_Y05_reset_out;
wire [0:0] Tile_X0A_Y05_stall_out;
wire [7:0] Tile_X0A_Y05_lo_out;
wire [15:0] Tile_X0A_Y05_tile_id_in;
wire [0:0] Tile_X0A_Y06_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y06_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y06_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y06_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y06_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y06_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y06_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y06_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y06_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y06_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y06_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y06_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y06_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y06_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y06_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y06_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y06_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y06_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y06_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y06_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y06_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y06_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y06_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y06_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y06_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y06_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y06_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y06_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y06_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y06_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y06_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y06_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y06_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y06_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y06_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y06_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y06_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y06_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y06_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y06_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0A_Y06_clk_out;
wire Tile_X0A_Y06_clk_pass_through_out_bot;
wire Tile_X0A_Y06_clk_pass_through_out_right;
wire [31:0] Tile_X0A_Y06_config_out_config_addr;
wire [31:0] Tile_X0A_Y06_config_out_config_data;
wire [0:0] Tile_X0A_Y06_config_out_read;
wire [0:0] Tile_X0A_Y06_config_out_write;
wire [8:0] Tile_X0A_Y06_hi;
wire [7:0] Tile_X0A_Y06_lo_unq1;
wire [31:0] Tile_X0A_Y06_read_config_data;
wire Tile_X0A_Y06_reset_out;
wire [0:0] Tile_X0A_Y06_stall_out;
wire [7:0] Tile_X0A_Y06_lo_out;
wire [15:0] Tile_X0A_Y06_tile_id_in;
wire [0:0] Tile_X0A_Y07_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y07_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y07_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y07_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y07_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y07_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y07_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y07_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y07_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y07_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y07_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y07_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y07_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y07_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y07_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y07_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y07_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y07_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y07_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y07_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y07_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y07_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y07_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y07_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y07_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y07_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y07_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y07_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y07_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y07_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y07_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y07_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y07_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y07_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y07_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y07_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y07_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y07_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y07_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y07_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0A_Y07_clk_out;
wire Tile_X0A_Y07_clk_pass_through_out_bot;
wire Tile_X0A_Y07_clk_pass_through_out_right;
wire [31:0] Tile_X0A_Y07_config_out_config_addr;
wire [31:0] Tile_X0A_Y07_config_out_config_data;
wire [0:0] Tile_X0A_Y07_config_out_read;
wire [0:0] Tile_X0A_Y07_config_out_write;
wire [8:0] Tile_X0A_Y07_hi_unq1;
wire [7:0] Tile_X0A_Y07_lo_unq1;
wire [31:0] Tile_X0A_Y07_read_config_data;
wire Tile_X0A_Y07_reset_out;
wire [0:0] Tile_X0A_Y07_stall_out;
wire [8:0] Tile_X0A_Y07_hi_out;
wire [7:0] Tile_X0A_Y07_lo_out;
wire [15:0] Tile_X0A_Y07_tile_id_in;
wire [0:0] Tile_X0A_Y08_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y08_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y08_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y08_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y08_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y08_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y08_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y08_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y08_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y08_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y08_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y08_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y08_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y08_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y08_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y08_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y08_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y08_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y08_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y08_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y08_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y08_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y08_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y08_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y08_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y08_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y08_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y08_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y08_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y08_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y08_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y08_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y08_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y08_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y08_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y08_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y08_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y08_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y08_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y08_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0A_Y08_clk_out;
wire Tile_X0A_Y08_clk_pass_through_out_bot;
wire Tile_X0A_Y08_clk_pass_through_out_right;
wire [31:0] Tile_X0A_Y08_config_out_config_addr;
wire [31:0] Tile_X0A_Y08_config_out_config_data;
wire [0:0] Tile_X0A_Y08_config_out_read;
wire [0:0] Tile_X0A_Y08_config_out_write;
wire [8:0] Tile_X0A_Y08_hi;
wire [7:0] Tile_X0A_Y08_lo_unq1;
wire [31:0] Tile_X0A_Y08_read_config_data;
wire Tile_X0A_Y08_reset_out;
wire [0:0] Tile_X0A_Y08_stall_out;
wire [7:0] Tile_X0A_Y08_lo_out;
wire [15:0] Tile_X0A_Y08_tile_id_in;
wire [0:0] Tile_X0A_Y09_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y09_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y09_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y09_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y09_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y09_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y09_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y09_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y09_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y09_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y09_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y09_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y09_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y09_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y09_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y09_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y09_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y09_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y09_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y09_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y09_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y09_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y09_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y09_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y09_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y09_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y09_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y09_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y09_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y09_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y09_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y09_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y09_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y09_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y09_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y09_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y09_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y09_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y09_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y09_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0A_Y09_clk_out;
wire Tile_X0A_Y09_clk_pass_through_out_bot;
wire Tile_X0A_Y09_clk_pass_through_out_right;
wire [31:0] Tile_X0A_Y09_config_out_config_addr;
wire [31:0] Tile_X0A_Y09_config_out_config_data;
wire [0:0] Tile_X0A_Y09_config_out_read;
wire [0:0] Tile_X0A_Y09_config_out_write;
wire [8:0] Tile_X0A_Y09_hi;
wire [7:0] Tile_X0A_Y09_lo_unq1;
wire [31:0] Tile_X0A_Y09_read_config_data;
wire Tile_X0A_Y09_reset_out;
wire [0:0] Tile_X0A_Y09_stall_out;
wire [7:0] Tile_X0A_Y09_lo_out;
wire [15:0] Tile_X0A_Y09_tile_id_in;
wire [0:0] Tile_X0A_Y0A_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0A_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0A_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0A_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0A_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0A_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0A_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0A_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0A_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0A_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0A_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0A_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0A_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0A_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0A_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0A_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0A_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0A_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0A_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0A_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0A_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0A_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0A_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0A_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0A_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0A_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0A_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0A_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0A_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0A_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0A_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0A_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0A_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0A_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0A_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0A_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0A_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0A_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0A_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0A_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0A_Y0A_clk_out;
wire Tile_X0A_Y0A_clk_pass_through_out_bot;
wire Tile_X0A_Y0A_clk_pass_through_out_right;
wire [31:0] Tile_X0A_Y0A_config_out_config_addr;
wire [31:0] Tile_X0A_Y0A_config_out_config_data;
wire [0:0] Tile_X0A_Y0A_config_out_read;
wire [0:0] Tile_X0A_Y0A_config_out_write;
wire [8:0] Tile_X0A_Y0A_hi;
wire [7:0] Tile_X0A_Y0A_lo_unq1;
wire [31:0] Tile_X0A_Y0A_read_config_data;
wire Tile_X0A_Y0A_reset_out;
wire [0:0] Tile_X0A_Y0A_stall_out;
wire [7:0] Tile_X0A_Y0A_lo_out;
wire [15:0] Tile_X0A_Y0A_tile_id_in;
wire [0:0] Tile_X0A_Y0B_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0B_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0B_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0B_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0B_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0B_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0B_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0B_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0B_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0B_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0B_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0B_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0B_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0B_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0B_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0B_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0B_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0B_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0B_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0B_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0B_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0B_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0B_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0B_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0B_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0B_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0B_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0B_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0B_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0B_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0B_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0B_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0B_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0B_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0B_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0B_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0B_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0B_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0B_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0B_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0A_Y0B_clk_out;
wire Tile_X0A_Y0B_clk_pass_through_out_bot;
wire Tile_X0A_Y0B_clk_pass_through_out_right;
wire [31:0] Tile_X0A_Y0B_config_out_config_addr;
wire [31:0] Tile_X0A_Y0B_config_out_config_data;
wire [0:0] Tile_X0A_Y0B_config_out_read;
wire [0:0] Tile_X0A_Y0B_config_out_write;
wire [8:0] Tile_X0A_Y0B_hi_unq1;
wire [7:0] Tile_X0A_Y0B_lo_unq1;
wire [31:0] Tile_X0A_Y0B_read_config_data;
wire Tile_X0A_Y0B_reset_out;
wire [0:0] Tile_X0A_Y0B_stall_out;
wire [8:0] Tile_X0A_Y0B_hi_out;
wire [7:0] Tile_X0A_Y0B_lo_out;
wire [15:0] Tile_X0A_Y0B_tile_id_in;
wire [0:0] Tile_X0A_Y0C_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0C_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0C_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0C_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0C_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0C_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0C_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0C_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0C_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0C_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0C_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0C_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0C_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0C_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0C_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0C_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0C_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0C_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0C_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0C_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0C_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0C_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0C_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0C_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0C_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0C_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0C_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0C_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0C_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0C_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0C_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0C_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0C_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0C_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0C_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0C_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0C_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0C_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0C_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0C_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0A_Y0C_clk_out;
wire Tile_X0A_Y0C_clk_pass_through_out_bot;
wire Tile_X0A_Y0C_clk_pass_through_out_right;
wire [31:0] Tile_X0A_Y0C_config_out_config_addr;
wire [31:0] Tile_X0A_Y0C_config_out_config_data;
wire [0:0] Tile_X0A_Y0C_config_out_read;
wire [0:0] Tile_X0A_Y0C_config_out_write;
wire [8:0] Tile_X0A_Y0C_hi_unq1;
wire [7:0] Tile_X0A_Y0C_lo_unq1;
wire [31:0] Tile_X0A_Y0C_read_config_data;
wire Tile_X0A_Y0C_reset_out;
wire [0:0] Tile_X0A_Y0C_stall_out;
wire [8:0] Tile_X0A_Y0C_hi_out;
wire [7:0] Tile_X0A_Y0C_lo_out;
wire [15:0] Tile_X0A_Y0C_tile_id_in;
wire [0:0] Tile_X0A_Y0D_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0D_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0D_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0D_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0D_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0D_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0D_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0D_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0D_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0D_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0D_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0D_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0D_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0D_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0D_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0D_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0D_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0D_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0D_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0D_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0D_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0D_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0D_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0D_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0D_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0D_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0D_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0D_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0D_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0D_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0D_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0D_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0D_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0D_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0D_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0D_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0D_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0D_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0D_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0D_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0A_Y0D_clk_out;
wire Tile_X0A_Y0D_clk_pass_through_out_bot;
wire Tile_X0A_Y0D_clk_pass_through_out_right;
wire [31:0] Tile_X0A_Y0D_config_out_config_addr;
wire [31:0] Tile_X0A_Y0D_config_out_config_data;
wire [0:0] Tile_X0A_Y0D_config_out_read;
wire [0:0] Tile_X0A_Y0D_config_out_write;
wire [8:0] Tile_X0A_Y0D_hi_unq1;
wire [7:0] Tile_X0A_Y0D_lo_unq1;
wire [31:0] Tile_X0A_Y0D_read_config_data;
wire Tile_X0A_Y0D_reset_out;
wire [0:0] Tile_X0A_Y0D_stall_out;
wire [8:0] Tile_X0A_Y0D_hi_out;
wire [7:0] Tile_X0A_Y0D_lo_out;
wire [15:0] Tile_X0A_Y0D_tile_id_in;
wire [0:0] Tile_X0A_Y0E_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0E_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0E_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0E_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0E_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0E_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0E_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0E_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0E_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0E_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0E_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0E_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0E_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0E_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0E_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0E_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0E_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0E_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0E_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0E_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0E_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0E_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0E_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0E_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0E_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0E_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0E_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0E_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0E_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0E_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0E_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0E_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0E_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0E_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0E_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0E_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0E_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0E_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0E_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0E_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0A_Y0E_clk_out;
wire Tile_X0A_Y0E_clk_pass_through_out_bot;
wire Tile_X0A_Y0E_clk_pass_through_out_right;
wire [31:0] Tile_X0A_Y0E_config_out_config_addr;
wire [31:0] Tile_X0A_Y0E_config_out_config_data;
wire [0:0] Tile_X0A_Y0E_config_out_read;
wire [0:0] Tile_X0A_Y0E_config_out_write;
wire [8:0] Tile_X0A_Y0E_hi_unq1;
wire [7:0] Tile_X0A_Y0E_lo_unq1;
wire [31:0] Tile_X0A_Y0E_read_config_data;
wire Tile_X0A_Y0E_reset_out;
wire [0:0] Tile_X0A_Y0E_stall_out;
wire [8:0] Tile_X0A_Y0E_hi_out;
wire [7:0] Tile_X0A_Y0E_lo_out;
wire [15:0] Tile_X0A_Y0E_tile_id_in;
wire [0:0] Tile_X0A_Y0F_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0F_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0F_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0F_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0F_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0F_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0F_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0F_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0F_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0F_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0F_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0F_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0F_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0F_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0F_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0F_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0F_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0F_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0F_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0F_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0F_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0F_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0F_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0F_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0F_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0F_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0F_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0F_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0F_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0F_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0F_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0F_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0F_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0F_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0F_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0F_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0F_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0F_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y0F_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y0F_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0A_Y0F_clk_out;
wire Tile_X0A_Y0F_clk_pass_through_out_bot;
wire Tile_X0A_Y0F_clk_pass_through_out_right;
wire [31:0] Tile_X0A_Y0F_config_out_config_addr;
wire [31:0] Tile_X0A_Y0F_config_out_config_data;
wire [0:0] Tile_X0A_Y0F_config_out_read;
wire [0:0] Tile_X0A_Y0F_config_out_write;
wire [8:0] Tile_X0A_Y0F_hi_unq1;
wire [7:0] Tile_X0A_Y0F_lo_unq1;
wire [31:0] Tile_X0A_Y0F_read_config_data;
wire Tile_X0A_Y0F_reset_out;
wire [0:0] Tile_X0A_Y0F_stall_out;
wire [8:0] Tile_X0A_Y0F_hi_out;
wire [7:0] Tile_X0A_Y0F_lo_out;
wire [15:0] Tile_X0A_Y0F_tile_id_in;
wire [0:0] Tile_X0A_Y10_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y10_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y10_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y10_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y10_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y10_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y10_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y10_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y10_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y10_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y10_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y10_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y10_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y10_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y10_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y10_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y10_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y10_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y10_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y10_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y10_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y10_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y10_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y10_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y10_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y10_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y10_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y10_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y10_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y10_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y10_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y10_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y10_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y10_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0A_Y10_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y10_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y10_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0A_Y10_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0A_Y10_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0A_Y10_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0A_Y10_clk_out;
wire Tile_X0A_Y10_clk_pass_through_out_bot;
wire Tile_X0A_Y10_clk_pass_through_out_right;
wire [31:0] Tile_X0A_Y10_config_out_config_addr;
wire [31:0] Tile_X0A_Y10_config_out_config_data;
wire [0:0] Tile_X0A_Y10_config_out_read;
wire [0:0] Tile_X0A_Y10_config_out_write;
wire [8:0] Tile_X0A_Y10_hi;
wire [7:0] Tile_X0A_Y10_lo_unq1;
wire [31:0] Tile_X0A_Y10_read_config_data;
wire Tile_X0A_Y10_reset_out;
wire [0:0] Tile_X0A_Y10_stall_out;
wire [7:0] Tile_X0A_Y10_lo_out;
wire [15:0] Tile_X0A_Y10_tile_id_in;
wire [0:0] Tile_X0B_Y00_io2glb_1;
wire [0:0] Tile_X0B_Y00_io2f_1;
wire [15:0] Tile_X0B_Y00_io2glb_16;
wire [15:0] Tile_X0B_Y00_io2f_16;
wire [8:0] Tile_X0B_Y00_hi;
wire [7:0] Tile_X0B_Y00_lo;
wire [0:0] Tile_X0B_Y01_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y01_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y01_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y01_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y01_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y01_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y01_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y01_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y01_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y01_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y01_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y01_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y01_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y01_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y01_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y01_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y01_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y01_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y01_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y01_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y01_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y01_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y01_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y01_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y01_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y01_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y01_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y01_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y01_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y01_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y01_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y01_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y01_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y01_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y01_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y01_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y01_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y01_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y01_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y01_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0B_Y01_clk_out;
wire [31:0] Tile_X0B_Y01_config_out_config_addr;
wire [31:0] Tile_X0B_Y01_config_out_config_data;
wire [0:0] Tile_X0B_Y01_config_out_read;
wire [0:0] Tile_X0B_Y01_config_out_write;
wire [8:0] Tile_X0B_Y01_hi_unq1;
wire [7:0] Tile_X0B_Y01_lo_unq1;
wire [31:0] Tile_X0B_Y01_read_config_data;
wire Tile_X0B_Y01_reset_out;
wire [0:0] Tile_X0B_Y01_stall_out;
wire [8:0] Tile_X0B_Y01_hi_out;
wire [7:0] Tile_X0B_Y01_lo_out;
wire [15:0] Tile_X0B_Y01_tile_id_in;
wire [0:0] Tile_X0B_Y02_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y02_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y02_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y02_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y02_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y02_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y02_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y02_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y02_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y02_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y02_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y02_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y02_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y02_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y02_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y02_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y02_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y02_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y02_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y02_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y02_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y02_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y02_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y02_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y02_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y02_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y02_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y02_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y02_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y02_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y02_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y02_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y02_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y02_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y02_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y02_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y02_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y02_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y02_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y02_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0B_Y02_clk_out;
wire [31:0] Tile_X0B_Y02_config_out_config_addr;
wire [31:0] Tile_X0B_Y02_config_out_config_data;
wire [0:0] Tile_X0B_Y02_config_out_read;
wire [0:0] Tile_X0B_Y02_config_out_write;
wire [8:0] Tile_X0B_Y02_hi_unq1;
wire [7:0] Tile_X0B_Y02_lo_unq1;
wire [31:0] Tile_X0B_Y02_read_config_data;
wire Tile_X0B_Y02_reset_out;
wire [0:0] Tile_X0B_Y02_stall_out;
wire [8:0] Tile_X0B_Y02_hi_out;
wire [7:0] Tile_X0B_Y02_lo_out;
wire [15:0] Tile_X0B_Y02_tile_id_in;
wire [0:0] Tile_X0B_Y03_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y03_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y03_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y03_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y03_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y03_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y03_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y03_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y03_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y03_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y03_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y03_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y03_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y03_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y03_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y03_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y03_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y03_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y03_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y03_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y03_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y03_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y03_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y03_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y03_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y03_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y03_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y03_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y03_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y03_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y03_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y03_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y03_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y03_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y03_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y03_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y03_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y03_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y03_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y03_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0B_Y03_clk_out;
wire [31:0] Tile_X0B_Y03_config_out_config_addr;
wire [31:0] Tile_X0B_Y03_config_out_config_data;
wire [0:0] Tile_X0B_Y03_config_out_read;
wire [0:0] Tile_X0B_Y03_config_out_write;
wire [8:0] Tile_X0B_Y03_hi_unq1;
wire [7:0] Tile_X0B_Y03_lo_unq1;
wire [31:0] Tile_X0B_Y03_read_config_data;
wire Tile_X0B_Y03_reset_out;
wire [0:0] Tile_X0B_Y03_stall_out;
wire [8:0] Tile_X0B_Y03_hi_out;
wire [7:0] Tile_X0B_Y03_lo_out;
wire [15:0] Tile_X0B_Y03_tile_id_in;
wire [0:0] Tile_X0B_Y04_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y04_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y04_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y04_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y04_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y04_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y04_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y04_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y04_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y04_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y04_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y04_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y04_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y04_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y04_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y04_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y04_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y04_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y04_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y04_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y04_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y04_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y04_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y04_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y04_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y04_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y04_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y04_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y04_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y04_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y04_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y04_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y04_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y04_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y04_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y04_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y04_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y04_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y04_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y04_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0B_Y04_clk_out;
wire [31:0] Tile_X0B_Y04_config_out_config_addr;
wire [31:0] Tile_X0B_Y04_config_out_config_data;
wire [0:0] Tile_X0B_Y04_config_out_read;
wire [0:0] Tile_X0B_Y04_config_out_write;
wire [8:0] Tile_X0B_Y04_hi_unq1;
wire [7:0] Tile_X0B_Y04_lo_unq1;
wire [31:0] Tile_X0B_Y04_read_config_data;
wire Tile_X0B_Y04_reset_out;
wire [0:0] Tile_X0B_Y04_stall_out;
wire [8:0] Tile_X0B_Y04_hi_out;
wire [7:0] Tile_X0B_Y04_lo_out;
wire [15:0] Tile_X0B_Y04_tile_id_in;
wire [0:0] Tile_X0B_Y05_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y05_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y05_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y05_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y05_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y05_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y05_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y05_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y05_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y05_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y05_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y05_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y05_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y05_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y05_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y05_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y05_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y05_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y05_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y05_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y05_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y05_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y05_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y05_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y05_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y05_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y05_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y05_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y05_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y05_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y05_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y05_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y05_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y05_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y05_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y05_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y05_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y05_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y05_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y05_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0B_Y05_clk_out;
wire [31:0] Tile_X0B_Y05_config_out_config_addr;
wire [31:0] Tile_X0B_Y05_config_out_config_data;
wire [0:0] Tile_X0B_Y05_config_out_read;
wire [0:0] Tile_X0B_Y05_config_out_write;
wire [8:0] Tile_X0B_Y05_hi_unq1;
wire [7:0] Tile_X0B_Y05_lo_unq1;
wire [31:0] Tile_X0B_Y05_read_config_data;
wire Tile_X0B_Y05_reset_out;
wire [0:0] Tile_X0B_Y05_stall_out;
wire [8:0] Tile_X0B_Y05_hi_out;
wire [7:0] Tile_X0B_Y05_lo_out;
wire [15:0] Tile_X0B_Y05_tile_id_in;
wire [0:0] Tile_X0B_Y06_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y06_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y06_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y06_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y06_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y06_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y06_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y06_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y06_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y06_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y06_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y06_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y06_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y06_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y06_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y06_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y06_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y06_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y06_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y06_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y06_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y06_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y06_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y06_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y06_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y06_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y06_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y06_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y06_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y06_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y06_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y06_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y06_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y06_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y06_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y06_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y06_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y06_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y06_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y06_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0B_Y06_clk_out;
wire [31:0] Tile_X0B_Y06_config_out_config_addr;
wire [31:0] Tile_X0B_Y06_config_out_config_data;
wire [0:0] Tile_X0B_Y06_config_out_read;
wire [0:0] Tile_X0B_Y06_config_out_write;
wire [8:0] Tile_X0B_Y06_hi_unq1;
wire [7:0] Tile_X0B_Y06_lo_unq1;
wire [31:0] Tile_X0B_Y06_read_config_data;
wire Tile_X0B_Y06_reset_out;
wire [0:0] Tile_X0B_Y06_stall_out;
wire [8:0] Tile_X0B_Y06_hi_out;
wire [7:0] Tile_X0B_Y06_lo_out;
wire [15:0] Tile_X0B_Y06_tile_id_in;
wire [0:0] Tile_X0B_Y07_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y07_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y07_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y07_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y07_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y07_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y07_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y07_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y07_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y07_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y07_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y07_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y07_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y07_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y07_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y07_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y07_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y07_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y07_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y07_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y07_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y07_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y07_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y07_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y07_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y07_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y07_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y07_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y07_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y07_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y07_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y07_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y07_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y07_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y07_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y07_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y07_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y07_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y07_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y07_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0B_Y07_clk_out;
wire [31:0] Tile_X0B_Y07_config_out_config_addr;
wire [31:0] Tile_X0B_Y07_config_out_config_data;
wire [0:0] Tile_X0B_Y07_config_out_read;
wire [0:0] Tile_X0B_Y07_config_out_write;
wire [8:0] Tile_X0B_Y07_hi_unq1;
wire [7:0] Tile_X0B_Y07_lo_unq1;
wire [31:0] Tile_X0B_Y07_read_config_data;
wire Tile_X0B_Y07_reset_out;
wire [0:0] Tile_X0B_Y07_stall_out;
wire [8:0] Tile_X0B_Y07_hi_out;
wire [7:0] Tile_X0B_Y07_lo_out;
wire [15:0] Tile_X0B_Y07_tile_id_in;
wire [0:0] Tile_X0B_Y08_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y08_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y08_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y08_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y08_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y08_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y08_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y08_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y08_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y08_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y08_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y08_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y08_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y08_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y08_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y08_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y08_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y08_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y08_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y08_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y08_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y08_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y08_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y08_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y08_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y08_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y08_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y08_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y08_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y08_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y08_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y08_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y08_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y08_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y08_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y08_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y08_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y08_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y08_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y08_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0B_Y08_clk_out;
wire [31:0] Tile_X0B_Y08_config_out_config_addr;
wire [31:0] Tile_X0B_Y08_config_out_config_data;
wire [0:0] Tile_X0B_Y08_config_out_read;
wire [0:0] Tile_X0B_Y08_config_out_write;
wire [8:0] Tile_X0B_Y08_hi_unq1;
wire [7:0] Tile_X0B_Y08_lo_unq1;
wire [31:0] Tile_X0B_Y08_read_config_data;
wire Tile_X0B_Y08_reset_out;
wire [0:0] Tile_X0B_Y08_stall_out;
wire [8:0] Tile_X0B_Y08_hi_out;
wire [7:0] Tile_X0B_Y08_lo_out;
wire [15:0] Tile_X0B_Y08_tile_id_in;
wire [0:0] Tile_X0B_Y09_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y09_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y09_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y09_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y09_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y09_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y09_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y09_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y09_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y09_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y09_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y09_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y09_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y09_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y09_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y09_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y09_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y09_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y09_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y09_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y09_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y09_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y09_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y09_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y09_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y09_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y09_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y09_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y09_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y09_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y09_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y09_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y09_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y09_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y09_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y09_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y09_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y09_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y09_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y09_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0B_Y09_clk_out;
wire [31:0] Tile_X0B_Y09_config_out_config_addr;
wire [31:0] Tile_X0B_Y09_config_out_config_data;
wire [0:0] Tile_X0B_Y09_config_out_read;
wire [0:0] Tile_X0B_Y09_config_out_write;
wire [8:0] Tile_X0B_Y09_hi_unq1;
wire [7:0] Tile_X0B_Y09_lo_unq1;
wire [31:0] Tile_X0B_Y09_read_config_data;
wire Tile_X0B_Y09_reset_out;
wire [0:0] Tile_X0B_Y09_stall_out;
wire [8:0] Tile_X0B_Y09_hi_out;
wire [7:0] Tile_X0B_Y09_lo_out;
wire [15:0] Tile_X0B_Y09_tile_id_in;
wire [0:0] Tile_X0B_Y0A_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0A_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0A_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0A_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0A_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0A_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0A_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0A_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0A_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0A_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0A_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0A_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0A_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0A_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0A_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0A_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0A_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0A_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0A_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0A_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0A_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0A_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0A_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0A_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0A_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0A_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0A_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0A_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0A_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0A_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0A_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0A_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0A_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0A_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0A_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0A_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0A_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0A_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0A_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0A_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0B_Y0A_clk_out;
wire [31:0] Tile_X0B_Y0A_config_out_config_addr;
wire [31:0] Tile_X0B_Y0A_config_out_config_data;
wire [0:0] Tile_X0B_Y0A_config_out_read;
wire [0:0] Tile_X0B_Y0A_config_out_write;
wire [8:0] Tile_X0B_Y0A_hi_unq1;
wire [7:0] Tile_X0B_Y0A_lo_unq1;
wire [31:0] Tile_X0B_Y0A_read_config_data;
wire Tile_X0B_Y0A_reset_out;
wire [0:0] Tile_X0B_Y0A_stall_out;
wire [8:0] Tile_X0B_Y0A_hi_out;
wire [7:0] Tile_X0B_Y0A_lo_out;
wire [15:0] Tile_X0B_Y0A_tile_id_in;
wire [0:0] Tile_X0B_Y0B_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0B_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0B_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0B_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0B_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0B_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0B_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0B_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0B_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0B_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0B_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0B_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0B_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0B_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0B_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0B_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0B_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0B_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0B_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0B_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0B_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0B_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0B_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0B_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0B_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0B_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0B_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0B_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0B_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0B_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0B_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0B_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0B_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0B_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0B_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0B_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0B_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0B_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0B_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0B_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0B_Y0B_clk_out;
wire [31:0] Tile_X0B_Y0B_config_out_config_addr;
wire [31:0] Tile_X0B_Y0B_config_out_config_data;
wire [0:0] Tile_X0B_Y0B_config_out_read;
wire [0:0] Tile_X0B_Y0B_config_out_write;
wire [8:0] Tile_X0B_Y0B_hi_unq1;
wire [7:0] Tile_X0B_Y0B_lo_unq1;
wire [31:0] Tile_X0B_Y0B_read_config_data;
wire Tile_X0B_Y0B_reset_out;
wire [0:0] Tile_X0B_Y0B_stall_out;
wire [8:0] Tile_X0B_Y0B_hi_out;
wire [7:0] Tile_X0B_Y0B_lo_out;
wire [15:0] Tile_X0B_Y0B_tile_id_in;
wire [0:0] Tile_X0B_Y0C_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0C_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0C_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0C_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0C_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0C_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0C_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0C_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0C_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0C_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0C_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0C_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0C_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0C_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0C_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0C_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0C_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0C_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0C_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0C_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0C_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0C_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0C_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0C_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0C_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0C_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0C_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0C_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0C_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0C_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0C_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0C_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0C_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0C_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0C_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0C_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0C_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0C_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0C_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0C_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0B_Y0C_clk_out;
wire [31:0] Tile_X0B_Y0C_config_out_config_addr;
wire [31:0] Tile_X0B_Y0C_config_out_config_data;
wire [0:0] Tile_X0B_Y0C_config_out_read;
wire [0:0] Tile_X0B_Y0C_config_out_write;
wire [8:0] Tile_X0B_Y0C_hi_unq1;
wire [7:0] Tile_X0B_Y0C_lo_unq1;
wire [31:0] Tile_X0B_Y0C_read_config_data;
wire Tile_X0B_Y0C_reset_out;
wire [0:0] Tile_X0B_Y0C_stall_out;
wire [8:0] Tile_X0B_Y0C_hi_out;
wire [7:0] Tile_X0B_Y0C_lo_out;
wire [15:0] Tile_X0B_Y0C_tile_id_in;
wire [0:0] Tile_X0B_Y0D_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0D_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0D_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0D_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0D_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0D_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0D_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0D_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0D_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0D_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0D_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0D_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0D_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0D_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0D_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0D_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0D_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0D_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0D_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0D_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0D_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0D_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0D_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0D_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0D_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0D_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0D_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0D_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0D_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0D_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0D_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0D_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0D_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0D_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0D_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0D_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0D_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0D_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0D_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0D_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0B_Y0D_clk_out;
wire [31:0] Tile_X0B_Y0D_config_out_config_addr;
wire [31:0] Tile_X0B_Y0D_config_out_config_data;
wire [0:0] Tile_X0B_Y0D_config_out_read;
wire [0:0] Tile_X0B_Y0D_config_out_write;
wire [8:0] Tile_X0B_Y0D_hi_unq1;
wire [7:0] Tile_X0B_Y0D_lo_unq1;
wire [31:0] Tile_X0B_Y0D_read_config_data;
wire Tile_X0B_Y0D_reset_out;
wire [0:0] Tile_X0B_Y0D_stall_out;
wire [8:0] Tile_X0B_Y0D_hi_out;
wire [7:0] Tile_X0B_Y0D_lo_out;
wire [15:0] Tile_X0B_Y0D_tile_id_in;
wire [0:0] Tile_X0B_Y0E_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0E_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0E_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0E_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0E_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0E_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0E_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0E_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0E_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0E_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0E_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0E_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0E_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0E_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0E_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0E_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0E_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0E_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0E_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0E_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0E_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0E_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0E_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0E_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0E_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0E_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0E_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0E_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0E_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0E_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0E_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0E_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0E_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0E_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0E_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0E_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0E_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0E_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0E_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0E_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0B_Y0E_clk_out;
wire [31:0] Tile_X0B_Y0E_config_out_config_addr;
wire [31:0] Tile_X0B_Y0E_config_out_config_data;
wire [0:0] Tile_X0B_Y0E_config_out_read;
wire [0:0] Tile_X0B_Y0E_config_out_write;
wire [8:0] Tile_X0B_Y0E_hi_unq1;
wire [7:0] Tile_X0B_Y0E_lo_unq1;
wire [31:0] Tile_X0B_Y0E_read_config_data;
wire Tile_X0B_Y0E_reset_out;
wire [0:0] Tile_X0B_Y0E_stall_out;
wire [8:0] Tile_X0B_Y0E_hi_out;
wire [7:0] Tile_X0B_Y0E_lo_out;
wire [15:0] Tile_X0B_Y0E_tile_id_in;
wire [0:0] Tile_X0B_Y0F_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0F_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0F_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0F_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0F_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0F_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0F_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0F_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0F_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0F_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0F_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0F_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0F_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0F_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0F_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0F_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0F_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0F_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0F_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0F_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0F_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0F_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0F_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0F_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0F_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0F_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0F_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0F_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0F_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0F_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0F_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0F_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0F_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0F_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0F_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0F_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0F_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0F_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y0F_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y0F_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0B_Y0F_clk_out;
wire [31:0] Tile_X0B_Y0F_config_out_config_addr;
wire [31:0] Tile_X0B_Y0F_config_out_config_data;
wire [0:0] Tile_X0B_Y0F_config_out_read;
wire [0:0] Tile_X0B_Y0F_config_out_write;
wire [8:0] Tile_X0B_Y0F_hi_unq1;
wire [7:0] Tile_X0B_Y0F_lo_unq1;
wire [31:0] Tile_X0B_Y0F_read_config_data;
wire Tile_X0B_Y0F_reset_out;
wire [0:0] Tile_X0B_Y0F_stall_out;
wire [8:0] Tile_X0B_Y0F_hi_out;
wire [7:0] Tile_X0B_Y0F_lo_out;
wire [15:0] Tile_X0B_Y0F_tile_id_in;
wire [0:0] Tile_X0B_Y10_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y10_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y10_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y10_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y10_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y10_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y10_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y10_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y10_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y10_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y10_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y10_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y10_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y10_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y10_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y10_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y10_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y10_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y10_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y10_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y10_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y10_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y10_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y10_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y10_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y10_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y10_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y10_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y10_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y10_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y10_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y10_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y10_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y10_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0B_Y10_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y10_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y10_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0B_Y10_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0B_Y10_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0B_Y10_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0B_Y10_clk_out;
wire [31:0] Tile_X0B_Y10_config_out_config_addr;
wire [31:0] Tile_X0B_Y10_config_out_config_data;
wire [0:0] Tile_X0B_Y10_config_out_read;
wire [0:0] Tile_X0B_Y10_config_out_write;
wire [8:0] Tile_X0B_Y10_hi_unq1;
wire [7:0] Tile_X0B_Y10_lo_unq1;
wire [31:0] Tile_X0B_Y10_read_config_data;
wire Tile_X0B_Y10_reset_out;
wire [0:0] Tile_X0B_Y10_stall_out;
wire [8:0] Tile_X0B_Y10_hi_out;
wire [7:0] Tile_X0B_Y10_lo_out;
wire [15:0] Tile_X0B_Y10_tile_id_in;
wire [0:0] Tile_X0C_Y00_io2glb_1;
wire [0:0] Tile_X0C_Y00_io2f_1;
wire [15:0] Tile_X0C_Y00_io2glb_16;
wire [15:0] Tile_X0C_Y00_io2f_16;
wire [8:0] Tile_X0C_Y00_hi;
wire [7:0] Tile_X0C_Y00_lo;
wire [0:0] Tile_X0C_Y01_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y01_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y01_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y01_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y01_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y01_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y01_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y01_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y01_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y01_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y01_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y01_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y01_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y01_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y01_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y01_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y01_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y01_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y01_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y01_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y01_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y01_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y01_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y01_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y01_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y01_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y01_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y01_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y01_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y01_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y01_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y01_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y01_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y01_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y01_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y01_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y01_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y01_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y01_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y01_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0C_Y01_clk_out;
wire Tile_X0C_Y01_clk_pass_through_out_bot;
wire Tile_X0C_Y01_clk_pass_through_out_right;
wire [31:0] Tile_X0C_Y01_config_out_config_addr;
wire [31:0] Tile_X0C_Y01_config_out_config_data;
wire [0:0] Tile_X0C_Y01_config_out_read;
wire [0:0] Tile_X0C_Y01_config_out_write;
wire [8:0] Tile_X0C_Y01_hi_unq1;
wire [7:0] Tile_X0C_Y01_lo_unq1;
wire [31:0] Tile_X0C_Y01_read_config_data;
wire Tile_X0C_Y01_reset_out;
wire [0:0] Tile_X0C_Y01_stall_out;
wire [8:0] Tile_X0C_Y01_hi_out;
wire [7:0] Tile_X0C_Y01_lo_out;
wire [15:0] Tile_X0C_Y01_tile_id_in;
wire [0:0] Tile_X0C_Y02_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y02_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y02_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y02_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y02_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y02_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y02_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y02_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y02_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y02_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y02_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y02_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y02_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y02_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y02_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y02_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y02_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y02_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y02_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y02_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y02_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y02_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y02_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y02_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y02_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y02_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y02_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y02_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y02_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y02_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y02_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y02_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y02_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y02_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y02_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y02_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y02_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y02_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y02_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y02_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0C_Y02_clk_out;
wire Tile_X0C_Y02_clk_pass_through_out_bot;
wire Tile_X0C_Y02_clk_pass_through_out_right;
wire [31:0] Tile_X0C_Y02_config_out_config_addr;
wire [31:0] Tile_X0C_Y02_config_out_config_data;
wire [0:0] Tile_X0C_Y02_config_out_read;
wire [0:0] Tile_X0C_Y02_config_out_write;
wire [8:0] Tile_X0C_Y02_hi_unq1;
wire [7:0] Tile_X0C_Y02_lo_unq1;
wire [31:0] Tile_X0C_Y02_read_config_data;
wire Tile_X0C_Y02_reset_out;
wire [0:0] Tile_X0C_Y02_stall_out;
wire [8:0] Tile_X0C_Y02_hi_out;
wire [7:0] Tile_X0C_Y02_lo_out;
wire [15:0] Tile_X0C_Y02_tile_id_in;
wire [0:0] Tile_X0C_Y03_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y03_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y03_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y03_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y03_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y03_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y03_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y03_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y03_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y03_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y03_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y03_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y03_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y03_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y03_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y03_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y03_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y03_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y03_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y03_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y03_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y03_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y03_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y03_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y03_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y03_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y03_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y03_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y03_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y03_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y03_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y03_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y03_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y03_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y03_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y03_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y03_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y03_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y03_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y03_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0C_Y03_clk_out;
wire Tile_X0C_Y03_clk_pass_through_out_bot;
wire Tile_X0C_Y03_clk_pass_through_out_right;
wire [31:0] Tile_X0C_Y03_config_out_config_addr;
wire [31:0] Tile_X0C_Y03_config_out_config_data;
wire [0:0] Tile_X0C_Y03_config_out_read;
wire [0:0] Tile_X0C_Y03_config_out_write;
wire [8:0] Tile_X0C_Y03_hi_unq1;
wire [7:0] Tile_X0C_Y03_lo_unq1;
wire [31:0] Tile_X0C_Y03_read_config_data;
wire Tile_X0C_Y03_reset_out;
wire [0:0] Tile_X0C_Y03_stall_out;
wire [8:0] Tile_X0C_Y03_hi_out;
wire [7:0] Tile_X0C_Y03_lo_out;
wire [15:0] Tile_X0C_Y03_tile_id_in;
wire [0:0] Tile_X0C_Y04_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y04_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y04_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y04_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y04_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y04_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y04_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y04_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y04_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y04_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y04_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y04_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y04_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y04_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y04_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y04_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y04_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y04_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y04_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y04_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y04_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y04_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y04_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y04_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y04_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y04_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y04_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y04_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y04_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y04_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y04_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y04_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y04_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y04_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y04_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y04_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y04_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y04_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y04_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y04_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0C_Y04_clk_out;
wire Tile_X0C_Y04_clk_pass_through_out_bot;
wire Tile_X0C_Y04_clk_pass_through_out_right;
wire [31:0] Tile_X0C_Y04_config_out_config_addr;
wire [31:0] Tile_X0C_Y04_config_out_config_data;
wire [0:0] Tile_X0C_Y04_config_out_read;
wire [0:0] Tile_X0C_Y04_config_out_write;
wire [8:0] Tile_X0C_Y04_hi_unq1;
wire [7:0] Tile_X0C_Y04_lo_unq1;
wire [31:0] Tile_X0C_Y04_read_config_data;
wire Tile_X0C_Y04_reset_out;
wire [0:0] Tile_X0C_Y04_stall_out;
wire [8:0] Tile_X0C_Y04_hi_out;
wire [7:0] Tile_X0C_Y04_lo_out;
wire [15:0] Tile_X0C_Y04_tile_id_in;
wire [0:0] Tile_X0C_Y05_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y05_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y05_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y05_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y05_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y05_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y05_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y05_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y05_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y05_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y05_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y05_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y05_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y05_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y05_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y05_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y05_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y05_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y05_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y05_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y05_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y05_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y05_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y05_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y05_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y05_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y05_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y05_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y05_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y05_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y05_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y05_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y05_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y05_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y05_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y05_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y05_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y05_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y05_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y05_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0C_Y05_clk_out;
wire Tile_X0C_Y05_clk_pass_through_out_bot;
wire Tile_X0C_Y05_clk_pass_through_out_right;
wire [31:0] Tile_X0C_Y05_config_out_config_addr;
wire [31:0] Tile_X0C_Y05_config_out_config_data;
wire [0:0] Tile_X0C_Y05_config_out_read;
wire [0:0] Tile_X0C_Y05_config_out_write;
wire [8:0] Tile_X0C_Y05_hi_unq1;
wire [7:0] Tile_X0C_Y05_lo_unq1;
wire [31:0] Tile_X0C_Y05_read_config_data;
wire Tile_X0C_Y05_reset_out;
wire [0:0] Tile_X0C_Y05_stall_out;
wire [8:0] Tile_X0C_Y05_hi_out;
wire [7:0] Tile_X0C_Y05_lo_out;
wire [15:0] Tile_X0C_Y05_tile_id_in;
wire [0:0] Tile_X0C_Y06_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y06_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y06_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y06_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y06_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y06_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y06_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y06_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y06_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y06_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y06_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y06_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y06_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y06_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y06_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y06_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y06_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y06_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y06_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y06_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y06_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y06_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y06_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y06_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y06_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y06_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y06_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y06_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y06_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y06_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y06_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y06_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y06_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y06_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y06_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y06_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y06_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y06_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y06_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y06_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0C_Y06_clk_out;
wire Tile_X0C_Y06_clk_pass_through_out_bot;
wire Tile_X0C_Y06_clk_pass_through_out_right;
wire [31:0] Tile_X0C_Y06_config_out_config_addr;
wire [31:0] Tile_X0C_Y06_config_out_config_data;
wire [0:0] Tile_X0C_Y06_config_out_read;
wire [0:0] Tile_X0C_Y06_config_out_write;
wire [8:0] Tile_X0C_Y06_hi_unq1;
wire [7:0] Tile_X0C_Y06_lo_unq1;
wire [31:0] Tile_X0C_Y06_read_config_data;
wire Tile_X0C_Y06_reset_out;
wire [0:0] Tile_X0C_Y06_stall_out;
wire [8:0] Tile_X0C_Y06_hi_out;
wire [7:0] Tile_X0C_Y06_lo_out;
wire [15:0] Tile_X0C_Y06_tile_id_in;
wire [0:0] Tile_X0C_Y07_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y07_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y07_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y07_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y07_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y07_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y07_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y07_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y07_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y07_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y07_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y07_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y07_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y07_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y07_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y07_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y07_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y07_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y07_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y07_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y07_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y07_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y07_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y07_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y07_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y07_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y07_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y07_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y07_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y07_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y07_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y07_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y07_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y07_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y07_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y07_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y07_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y07_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y07_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y07_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0C_Y07_clk_out;
wire Tile_X0C_Y07_clk_pass_through_out_bot;
wire Tile_X0C_Y07_clk_pass_through_out_right;
wire [31:0] Tile_X0C_Y07_config_out_config_addr;
wire [31:0] Tile_X0C_Y07_config_out_config_data;
wire [0:0] Tile_X0C_Y07_config_out_read;
wire [0:0] Tile_X0C_Y07_config_out_write;
wire [8:0] Tile_X0C_Y07_hi_unq1;
wire [7:0] Tile_X0C_Y07_lo_unq1;
wire [31:0] Tile_X0C_Y07_read_config_data;
wire Tile_X0C_Y07_reset_out;
wire [0:0] Tile_X0C_Y07_stall_out;
wire [8:0] Tile_X0C_Y07_hi_out;
wire [7:0] Tile_X0C_Y07_lo_out;
wire [15:0] Tile_X0C_Y07_tile_id_in;
wire [0:0] Tile_X0C_Y08_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y08_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y08_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y08_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y08_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y08_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y08_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y08_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y08_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y08_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y08_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y08_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y08_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y08_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y08_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y08_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y08_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y08_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y08_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y08_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y08_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y08_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y08_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y08_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y08_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y08_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y08_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y08_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y08_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y08_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y08_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y08_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y08_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y08_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y08_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y08_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y08_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y08_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y08_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y08_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0C_Y08_clk_out;
wire Tile_X0C_Y08_clk_pass_through_out_bot;
wire Tile_X0C_Y08_clk_pass_through_out_right;
wire [31:0] Tile_X0C_Y08_config_out_config_addr;
wire [31:0] Tile_X0C_Y08_config_out_config_data;
wire [0:0] Tile_X0C_Y08_config_out_read;
wire [0:0] Tile_X0C_Y08_config_out_write;
wire [8:0] Tile_X0C_Y08_hi_unq1;
wire [7:0] Tile_X0C_Y08_lo_unq1;
wire [31:0] Tile_X0C_Y08_read_config_data;
wire Tile_X0C_Y08_reset_out;
wire [0:0] Tile_X0C_Y08_stall_out;
wire [8:0] Tile_X0C_Y08_hi_out;
wire [7:0] Tile_X0C_Y08_lo_out;
wire [15:0] Tile_X0C_Y08_tile_id_in;
wire [0:0] Tile_X0C_Y09_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y09_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y09_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y09_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y09_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y09_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y09_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y09_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y09_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y09_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y09_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y09_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y09_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y09_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y09_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y09_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y09_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y09_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y09_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y09_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y09_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y09_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y09_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y09_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y09_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y09_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y09_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y09_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y09_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y09_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y09_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y09_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y09_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y09_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y09_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y09_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y09_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y09_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y09_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y09_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0C_Y09_clk_out;
wire Tile_X0C_Y09_clk_pass_through_out_bot;
wire Tile_X0C_Y09_clk_pass_through_out_right;
wire [31:0] Tile_X0C_Y09_config_out_config_addr;
wire [31:0] Tile_X0C_Y09_config_out_config_data;
wire [0:0] Tile_X0C_Y09_config_out_read;
wire [0:0] Tile_X0C_Y09_config_out_write;
wire [8:0] Tile_X0C_Y09_hi_unq1;
wire [7:0] Tile_X0C_Y09_lo_unq1;
wire [31:0] Tile_X0C_Y09_read_config_data;
wire Tile_X0C_Y09_reset_out;
wire [0:0] Tile_X0C_Y09_stall_out;
wire [8:0] Tile_X0C_Y09_hi_out;
wire [7:0] Tile_X0C_Y09_lo_out;
wire [15:0] Tile_X0C_Y09_tile_id_in;
wire [0:0] Tile_X0C_Y0A_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0A_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0A_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0A_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0A_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0A_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0A_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0A_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0A_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0A_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0A_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0A_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0A_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0A_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0A_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0A_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0A_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0A_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0A_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0A_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0A_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0A_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0A_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0A_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0A_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0A_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0A_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0A_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0A_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0A_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0A_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0A_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0A_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0A_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0A_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0A_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0A_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0A_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0A_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0A_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0C_Y0A_clk_out;
wire Tile_X0C_Y0A_clk_pass_through_out_bot;
wire Tile_X0C_Y0A_clk_pass_through_out_right;
wire [31:0] Tile_X0C_Y0A_config_out_config_addr;
wire [31:0] Tile_X0C_Y0A_config_out_config_data;
wire [0:0] Tile_X0C_Y0A_config_out_read;
wire [0:0] Tile_X0C_Y0A_config_out_write;
wire [8:0] Tile_X0C_Y0A_hi_unq1;
wire [7:0] Tile_X0C_Y0A_lo_unq1;
wire [31:0] Tile_X0C_Y0A_read_config_data;
wire Tile_X0C_Y0A_reset_out;
wire [0:0] Tile_X0C_Y0A_stall_out;
wire [8:0] Tile_X0C_Y0A_hi_out;
wire [7:0] Tile_X0C_Y0A_lo_out;
wire [15:0] Tile_X0C_Y0A_tile_id_in;
wire [0:0] Tile_X0C_Y0B_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0B_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0B_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0B_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0B_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0B_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0B_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0B_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0B_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0B_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0B_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0B_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0B_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0B_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0B_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0B_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0B_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0B_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0B_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0B_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0B_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0B_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0B_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0B_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0B_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0B_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0B_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0B_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0B_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0B_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0B_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0B_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0B_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0B_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0B_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0B_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0B_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0B_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0B_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0B_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0C_Y0B_clk_out;
wire Tile_X0C_Y0B_clk_pass_through_out_bot;
wire Tile_X0C_Y0B_clk_pass_through_out_right;
wire [31:0] Tile_X0C_Y0B_config_out_config_addr;
wire [31:0] Tile_X0C_Y0B_config_out_config_data;
wire [0:0] Tile_X0C_Y0B_config_out_read;
wire [0:0] Tile_X0C_Y0B_config_out_write;
wire [8:0] Tile_X0C_Y0B_hi_unq1;
wire [7:0] Tile_X0C_Y0B_lo_unq1;
wire [31:0] Tile_X0C_Y0B_read_config_data;
wire Tile_X0C_Y0B_reset_out;
wire [0:0] Tile_X0C_Y0B_stall_out;
wire [8:0] Tile_X0C_Y0B_hi_out;
wire [7:0] Tile_X0C_Y0B_lo_out;
wire [15:0] Tile_X0C_Y0B_tile_id_in;
wire [0:0] Tile_X0C_Y0C_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0C_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0C_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0C_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0C_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0C_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0C_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0C_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0C_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0C_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0C_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0C_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0C_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0C_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0C_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0C_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0C_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0C_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0C_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0C_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0C_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0C_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0C_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0C_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0C_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0C_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0C_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0C_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0C_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0C_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0C_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0C_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0C_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0C_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0C_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0C_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0C_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0C_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0C_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0C_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0C_Y0C_clk_out;
wire Tile_X0C_Y0C_clk_pass_through_out_bot;
wire Tile_X0C_Y0C_clk_pass_through_out_right;
wire [31:0] Tile_X0C_Y0C_config_out_config_addr;
wire [31:0] Tile_X0C_Y0C_config_out_config_data;
wire [0:0] Tile_X0C_Y0C_config_out_read;
wire [0:0] Tile_X0C_Y0C_config_out_write;
wire [8:0] Tile_X0C_Y0C_hi_unq1;
wire [7:0] Tile_X0C_Y0C_lo_unq1;
wire [31:0] Tile_X0C_Y0C_read_config_data;
wire Tile_X0C_Y0C_reset_out;
wire [0:0] Tile_X0C_Y0C_stall_out;
wire [8:0] Tile_X0C_Y0C_hi_out;
wire [7:0] Tile_X0C_Y0C_lo_out;
wire [15:0] Tile_X0C_Y0C_tile_id_in;
wire [0:0] Tile_X0C_Y0D_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0D_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0D_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0D_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0D_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0D_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0D_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0D_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0D_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0D_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0D_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0D_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0D_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0D_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0D_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0D_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0D_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0D_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0D_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0D_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0D_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0D_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0D_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0D_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0D_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0D_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0D_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0D_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0D_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0D_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0D_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0D_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0D_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0D_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0D_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0D_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0D_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0D_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0D_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0D_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0C_Y0D_clk_out;
wire Tile_X0C_Y0D_clk_pass_through_out_bot;
wire Tile_X0C_Y0D_clk_pass_through_out_right;
wire [31:0] Tile_X0C_Y0D_config_out_config_addr;
wire [31:0] Tile_X0C_Y0D_config_out_config_data;
wire [0:0] Tile_X0C_Y0D_config_out_read;
wire [0:0] Tile_X0C_Y0D_config_out_write;
wire [8:0] Tile_X0C_Y0D_hi_unq1;
wire [7:0] Tile_X0C_Y0D_lo_unq1;
wire [31:0] Tile_X0C_Y0D_read_config_data;
wire Tile_X0C_Y0D_reset_out;
wire [0:0] Tile_X0C_Y0D_stall_out;
wire [8:0] Tile_X0C_Y0D_hi_out;
wire [7:0] Tile_X0C_Y0D_lo_out;
wire [15:0] Tile_X0C_Y0D_tile_id_in;
wire [0:0] Tile_X0C_Y0E_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0E_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0E_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0E_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0E_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0E_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0E_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0E_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0E_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0E_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0E_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0E_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0E_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0E_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0E_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0E_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0E_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0E_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0E_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0E_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0E_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0E_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0E_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0E_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0E_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0E_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0E_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0E_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0E_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0E_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0E_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0E_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0E_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0E_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0E_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0E_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0E_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0E_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0E_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0E_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0C_Y0E_clk_out;
wire Tile_X0C_Y0E_clk_pass_through_out_bot;
wire Tile_X0C_Y0E_clk_pass_through_out_right;
wire [31:0] Tile_X0C_Y0E_config_out_config_addr;
wire [31:0] Tile_X0C_Y0E_config_out_config_data;
wire [0:0] Tile_X0C_Y0E_config_out_read;
wire [0:0] Tile_X0C_Y0E_config_out_write;
wire [8:0] Tile_X0C_Y0E_hi_unq1;
wire [7:0] Tile_X0C_Y0E_lo_unq1;
wire [31:0] Tile_X0C_Y0E_read_config_data;
wire Tile_X0C_Y0E_reset_out;
wire [0:0] Tile_X0C_Y0E_stall_out;
wire [8:0] Tile_X0C_Y0E_hi_out;
wire [7:0] Tile_X0C_Y0E_lo_out;
wire [15:0] Tile_X0C_Y0E_tile_id_in;
wire [0:0] Tile_X0C_Y0F_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0F_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0F_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0F_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0F_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0F_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0F_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0F_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0F_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0F_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0F_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0F_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0F_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0F_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0F_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0F_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0F_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0F_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0F_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0F_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0F_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0F_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0F_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0F_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0F_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0F_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0F_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0F_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0F_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0F_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0F_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0F_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0F_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0F_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0F_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0F_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0F_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0F_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y0F_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y0F_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0C_Y0F_clk_out;
wire Tile_X0C_Y0F_clk_pass_through_out_bot;
wire Tile_X0C_Y0F_clk_pass_through_out_right;
wire [31:0] Tile_X0C_Y0F_config_out_config_addr;
wire [31:0] Tile_X0C_Y0F_config_out_config_data;
wire [0:0] Tile_X0C_Y0F_config_out_read;
wire [0:0] Tile_X0C_Y0F_config_out_write;
wire [8:0] Tile_X0C_Y0F_hi_unq1;
wire [7:0] Tile_X0C_Y0F_lo_unq1;
wire [31:0] Tile_X0C_Y0F_read_config_data;
wire Tile_X0C_Y0F_reset_out;
wire [0:0] Tile_X0C_Y0F_stall_out;
wire [8:0] Tile_X0C_Y0F_hi_out;
wire [7:0] Tile_X0C_Y0F_lo_out;
wire [15:0] Tile_X0C_Y0F_tile_id_in;
wire [0:0] Tile_X0C_Y10_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y10_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y10_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y10_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y10_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y10_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y10_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y10_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y10_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y10_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y10_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y10_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y10_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y10_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y10_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y10_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y10_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y10_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y10_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y10_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y10_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y10_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y10_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y10_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y10_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y10_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y10_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y10_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y10_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y10_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y10_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y10_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y10_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y10_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0C_Y10_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y10_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y10_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0C_Y10_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0C_Y10_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0C_Y10_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0C_Y10_clk_out;
wire Tile_X0C_Y10_clk_pass_through_out_bot;
wire Tile_X0C_Y10_clk_pass_through_out_right;
wire [31:0] Tile_X0C_Y10_config_out_config_addr;
wire [31:0] Tile_X0C_Y10_config_out_config_data;
wire [0:0] Tile_X0C_Y10_config_out_read;
wire [0:0] Tile_X0C_Y10_config_out_write;
wire [8:0] Tile_X0C_Y10_hi_unq1;
wire [7:0] Tile_X0C_Y10_lo_unq1;
wire [31:0] Tile_X0C_Y10_read_config_data;
wire Tile_X0C_Y10_reset_out;
wire [0:0] Tile_X0C_Y10_stall_out;
wire [8:0] Tile_X0C_Y10_hi_out;
wire [7:0] Tile_X0C_Y10_lo_out;
wire [15:0] Tile_X0C_Y10_tile_id_in;
wire [0:0] Tile_X0D_Y00_io2glb_1;
wire [0:0] Tile_X0D_Y00_io2f_1;
wire [15:0] Tile_X0D_Y00_io2glb_16;
wire [15:0] Tile_X0D_Y00_io2f_16;
wire [8:0] Tile_X0D_Y00_hi;
wire [7:0] Tile_X0D_Y00_lo;
wire [0:0] Tile_X0D_Y01_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y01_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y01_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y01_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y01_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y01_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y01_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y01_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y01_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y01_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y01_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y01_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y01_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y01_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y01_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y01_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y01_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y01_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y01_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y01_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y01_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y01_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y01_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y01_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y01_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y01_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y01_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y01_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y01_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y01_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y01_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y01_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y01_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y01_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y01_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y01_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y01_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y01_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y01_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y01_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0D_Y01_clk_out;
wire Tile_X0D_Y01_clk_pass_through_out_bot;
wire Tile_X0D_Y01_clk_pass_through_out_right;
wire [31:0] Tile_X0D_Y01_config_out_config_addr;
wire [31:0] Tile_X0D_Y01_config_out_config_data;
wire [0:0] Tile_X0D_Y01_config_out_read;
wire [0:0] Tile_X0D_Y01_config_out_write;
wire [8:0] Tile_X0D_Y01_hi_unq1;
wire [7:0] Tile_X0D_Y01_lo_unq1;
wire [31:0] Tile_X0D_Y01_read_config_data;
wire Tile_X0D_Y01_reset_out;
wire [0:0] Tile_X0D_Y01_stall_out;
wire [8:0] Tile_X0D_Y01_hi_out;
wire [7:0] Tile_X0D_Y01_lo_out;
wire [15:0] Tile_X0D_Y01_tile_id_in;
wire [0:0] Tile_X0D_Y02_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y02_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y02_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y02_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y02_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y02_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y02_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y02_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y02_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y02_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y02_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y02_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y02_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y02_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y02_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y02_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y02_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y02_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y02_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y02_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y02_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y02_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y02_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y02_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y02_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y02_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y02_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y02_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y02_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y02_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y02_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y02_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y02_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y02_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y02_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y02_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y02_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y02_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y02_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y02_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0D_Y02_clk_out;
wire Tile_X0D_Y02_clk_pass_through_out_bot;
wire Tile_X0D_Y02_clk_pass_through_out_right;
wire [31:0] Tile_X0D_Y02_config_out_config_addr;
wire [31:0] Tile_X0D_Y02_config_out_config_data;
wire [0:0] Tile_X0D_Y02_config_out_read;
wire [0:0] Tile_X0D_Y02_config_out_write;
wire [8:0] Tile_X0D_Y02_hi_unq1;
wire [7:0] Tile_X0D_Y02_lo_unq1;
wire [31:0] Tile_X0D_Y02_read_config_data;
wire Tile_X0D_Y02_reset_out;
wire [0:0] Tile_X0D_Y02_stall_out;
wire [8:0] Tile_X0D_Y02_hi_out;
wire [7:0] Tile_X0D_Y02_lo_out;
wire [15:0] Tile_X0D_Y02_tile_id_in;
wire [0:0] Tile_X0D_Y03_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y03_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y03_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y03_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y03_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y03_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y03_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y03_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y03_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y03_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y03_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y03_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y03_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y03_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y03_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y03_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y03_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y03_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y03_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y03_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y03_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y03_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y03_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y03_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y03_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y03_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y03_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y03_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y03_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y03_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y03_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y03_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y03_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y03_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y03_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y03_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y03_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y03_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y03_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y03_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0D_Y03_clk_out;
wire Tile_X0D_Y03_clk_pass_through_out_bot;
wire Tile_X0D_Y03_clk_pass_through_out_right;
wire [31:0] Tile_X0D_Y03_config_out_config_addr;
wire [31:0] Tile_X0D_Y03_config_out_config_data;
wire [0:0] Tile_X0D_Y03_config_out_read;
wire [0:0] Tile_X0D_Y03_config_out_write;
wire [8:0] Tile_X0D_Y03_hi_unq1;
wire [7:0] Tile_X0D_Y03_lo_unq1;
wire [31:0] Tile_X0D_Y03_read_config_data;
wire Tile_X0D_Y03_reset_out;
wire [0:0] Tile_X0D_Y03_stall_out;
wire [8:0] Tile_X0D_Y03_hi_out;
wire [7:0] Tile_X0D_Y03_lo_out;
wire [15:0] Tile_X0D_Y03_tile_id_in;
wire [0:0] Tile_X0D_Y04_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y04_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y04_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y04_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y04_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y04_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y04_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y04_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y04_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y04_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y04_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y04_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y04_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y04_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y04_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y04_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y04_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y04_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y04_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y04_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y04_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y04_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y04_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y04_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y04_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y04_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y04_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y04_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y04_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y04_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y04_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y04_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y04_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y04_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y04_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y04_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y04_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y04_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y04_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y04_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0D_Y04_clk_out;
wire Tile_X0D_Y04_clk_pass_through_out_bot;
wire Tile_X0D_Y04_clk_pass_through_out_right;
wire [31:0] Tile_X0D_Y04_config_out_config_addr;
wire [31:0] Tile_X0D_Y04_config_out_config_data;
wire [0:0] Tile_X0D_Y04_config_out_read;
wire [0:0] Tile_X0D_Y04_config_out_write;
wire [8:0] Tile_X0D_Y04_hi_unq1;
wire [7:0] Tile_X0D_Y04_lo_unq1;
wire [31:0] Tile_X0D_Y04_read_config_data;
wire Tile_X0D_Y04_reset_out;
wire [0:0] Tile_X0D_Y04_stall_out;
wire [8:0] Tile_X0D_Y04_hi_out;
wire [7:0] Tile_X0D_Y04_lo_out;
wire [15:0] Tile_X0D_Y04_tile_id_in;
wire [0:0] Tile_X0D_Y05_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y05_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y05_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y05_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y05_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y05_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y05_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y05_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y05_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y05_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y05_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y05_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y05_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y05_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y05_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y05_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y05_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y05_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y05_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y05_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y05_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y05_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y05_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y05_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y05_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y05_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y05_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y05_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y05_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y05_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y05_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y05_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y05_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y05_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y05_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y05_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y05_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y05_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y05_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y05_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0D_Y05_clk_out;
wire Tile_X0D_Y05_clk_pass_through_out_bot;
wire Tile_X0D_Y05_clk_pass_through_out_right;
wire [31:0] Tile_X0D_Y05_config_out_config_addr;
wire [31:0] Tile_X0D_Y05_config_out_config_data;
wire [0:0] Tile_X0D_Y05_config_out_read;
wire [0:0] Tile_X0D_Y05_config_out_write;
wire [8:0] Tile_X0D_Y05_hi_unq1;
wire [7:0] Tile_X0D_Y05_lo_unq1;
wire [31:0] Tile_X0D_Y05_read_config_data;
wire Tile_X0D_Y05_reset_out;
wire [0:0] Tile_X0D_Y05_stall_out;
wire [8:0] Tile_X0D_Y05_hi_out;
wire [7:0] Tile_X0D_Y05_lo_out;
wire [15:0] Tile_X0D_Y05_tile_id_in;
wire [0:0] Tile_X0D_Y06_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y06_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y06_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y06_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y06_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y06_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y06_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y06_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y06_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y06_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y06_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y06_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y06_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y06_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y06_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y06_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y06_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y06_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y06_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y06_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y06_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y06_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y06_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y06_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y06_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y06_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y06_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y06_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y06_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y06_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y06_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y06_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y06_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y06_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y06_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y06_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y06_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y06_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y06_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y06_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0D_Y06_clk_out;
wire Tile_X0D_Y06_clk_pass_through_out_bot;
wire Tile_X0D_Y06_clk_pass_through_out_right;
wire [31:0] Tile_X0D_Y06_config_out_config_addr;
wire [31:0] Tile_X0D_Y06_config_out_config_data;
wire [0:0] Tile_X0D_Y06_config_out_read;
wire [0:0] Tile_X0D_Y06_config_out_write;
wire [8:0] Tile_X0D_Y06_hi_unq1;
wire [7:0] Tile_X0D_Y06_lo_unq1;
wire [31:0] Tile_X0D_Y06_read_config_data;
wire Tile_X0D_Y06_reset_out;
wire [0:0] Tile_X0D_Y06_stall_out;
wire [8:0] Tile_X0D_Y06_hi_out;
wire [7:0] Tile_X0D_Y06_lo_out;
wire [15:0] Tile_X0D_Y06_tile_id_in;
wire [0:0] Tile_X0D_Y07_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y07_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y07_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y07_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y07_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y07_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y07_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y07_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y07_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y07_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y07_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y07_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y07_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y07_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y07_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y07_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y07_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y07_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y07_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y07_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y07_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y07_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y07_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y07_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y07_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y07_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y07_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y07_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y07_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y07_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y07_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y07_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y07_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y07_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y07_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y07_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y07_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y07_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y07_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y07_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0D_Y07_clk_out;
wire Tile_X0D_Y07_clk_pass_through_out_bot;
wire Tile_X0D_Y07_clk_pass_through_out_right;
wire [31:0] Tile_X0D_Y07_config_out_config_addr;
wire [31:0] Tile_X0D_Y07_config_out_config_data;
wire [0:0] Tile_X0D_Y07_config_out_read;
wire [0:0] Tile_X0D_Y07_config_out_write;
wire [8:0] Tile_X0D_Y07_hi_unq1;
wire [7:0] Tile_X0D_Y07_lo_unq1;
wire [31:0] Tile_X0D_Y07_read_config_data;
wire Tile_X0D_Y07_reset_out;
wire [0:0] Tile_X0D_Y07_stall_out;
wire [8:0] Tile_X0D_Y07_hi_out;
wire [7:0] Tile_X0D_Y07_lo_out;
wire [15:0] Tile_X0D_Y07_tile_id_in;
wire [0:0] Tile_X0D_Y08_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y08_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y08_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y08_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y08_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y08_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y08_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y08_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y08_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y08_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y08_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y08_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y08_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y08_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y08_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y08_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y08_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y08_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y08_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y08_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y08_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y08_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y08_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y08_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y08_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y08_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y08_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y08_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y08_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y08_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y08_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y08_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y08_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y08_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y08_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y08_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y08_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y08_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y08_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y08_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0D_Y08_clk_out;
wire Tile_X0D_Y08_clk_pass_through_out_bot;
wire Tile_X0D_Y08_clk_pass_through_out_right;
wire [31:0] Tile_X0D_Y08_config_out_config_addr;
wire [31:0] Tile_X0D_Y08_config_out_config_data;
wire [0:0] Tile_X0D_Y08_config_out_read;
wire [0:0] Tile_X0D_Y08_config_out_write;
wire [8:0] Tile_X0D_Y08_hi_unq1;
wire [7:0] Tile_X0D_Y08_lo_unq1;
wire [31:0] Tile_X0D_Y08_read_config_data;
wire Tile_X0D_Y08_reset_out;
wire [0:0] Tile_X0D_Y08_stall_out;
wire [8:0] Tile_X0D_Y08_hi_out;
wire [7:0] Tile_X0D_Y08_lo_out;
wire [15:0] Tile_X0D_Y08_tile_id_in;
wire [0:0] Tile_X0D_Y09_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y09_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y09_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y09_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y09_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y09_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y09_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y09_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y09_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y09_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y09_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y09_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y09_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y09_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y09_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y09_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y09_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y09_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y09_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y09_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y09_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y09_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y09_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y09_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y09_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y09_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y09_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y09_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y09_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y09_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y09_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y09_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y09_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y09_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y09_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y09_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y09_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y09_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y09_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y09_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0D_Y09_clk_out;
wire Tile_X0D_Y09_clk_pass_through_out_bot;
wire Tile_X0D_Y09_clk_pass_through_out_right;
wire [31:0] Tile_X0D_Y09_config_out_config_addr;
wire [31:0] Tile_X0D_Y09_config_out_config_data;
wire [0:0] Tile_X0D_Y09_config_out_read;
wire [0:0] Tile_X0D_Y09_config_out_write;
wire [8:0] Tile_X0D_Y09_hi_unq1;
wire [7:0] Tile_X0D_Y09_lo_unq1;
wire [31:0] Tile_X0D_Y09_read_config_data;
wire Tile_X0D_Y09_reset_out;
wire [0:0] Tile_X0D_Y09_stall_out;
wire [8:0] Tile_X0D_Y09_hi_out;
wire [7:0] Tile_X0D_Y09_lo_out;
wire [15:0] Tile_X0D_Y09_tile_id_in;
wire [0:0] Tile_X0D_Y0A_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0A_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0A_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0A_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0A_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0A_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0A_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0A_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0A_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0A_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0A_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0A_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0A_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0A_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0A_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0A_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0A_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0A_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0A_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0A_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0A_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0A_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0A_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0A_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0A_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0A_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0A_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0A_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0A_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0A_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0A_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0A_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0A_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0A_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0A_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0A_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0A_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0A_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0A_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0A_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0D_Y0A_clk_out;
wire Tile_X0D_Y0A_clk_pass_through_out_bot;
wire Tile_X0D_Y0A_clk_pass_through_out_right;
wire [31:0] Tile_X0D_Y0A_config_out_config_addr;
wire [31:0] Tile_X0D_Y0A_config_out_config_data;
wire [0:0] Tile_X0D_Y0A_config_out_read;
wire [0:0] Tile_X0D_Y0A_config_out_write;
wire [8:0] Tile_X0D_Y0A_hi_unq1;
wire [7:0] Tile_X0D_Y0A_lo_unq1;
wire [31:0] Tile_X0D_Y0A_read_config_data;
wire Tile_X0D_Y0A_reset_out;
wire [0:0] Tile_X0D_Y0A_stall_out;
wire [8:0] Tile_X0D_Y0A_hi_out;
wire [7:0] Tile_X0D_Y0A_lo_out;
wire [15:0] Tile_X0D_Y0A_tile_id_in;
wire [0:0] Tile_X0D_Y0B_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0B_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0B_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0B_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0B_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0B_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0B_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0B_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0B_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0B_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0B_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0B_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0B_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0B_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0B_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0B_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0B_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0B_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0B_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0B_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0B_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0B_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0B_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0B_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0B_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0B_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0B_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0B_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0B_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0B_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0B_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0B_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0B_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0B_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0B_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0B_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0B_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0B_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0B_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0B_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0D_Y0B_clk_out;
wire Tile_X0D_Y0B_clk_pass_through_out_bot;
wire Tile_X0D_Y0B_clk_pass_through_out_right;
wire [31:0] Tile_X0D_Y0B_config_out_config_addr;
wire [31:0] Tile_X0D_Y0B_config_out_config_data;
wire [0:0] Tile_X0D_Y0B_config_out_read;
wire [0:0] Tile_X0D_Y0B_config_out_write;
wire [8:0] Tile_X0D_Y0B_hi_unq1;
wire [7:0] Tile_X0D_Y0B_lo_unq1;
wire [31:0] Tile_X0D_Y0B_read_config_data;
wire Tile_X0D_Y0B_reset_out;
wire [0:0] Tile_X0D_Y0B_stall_out;
wire [8:0] Tile_X0D_Y0B_hi_out;
wire [7:0] Tile_X0D_Y0B_lo_out;
wire [15:0] Tile_X0D_Y0B_tile_id_in;
wire [0:0] Tile_X0D_Y0C_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0C_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0C_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0C_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0C_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0C_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0C_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0C_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0C_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0C_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0C_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0C_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0C_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0C_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0C_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0C_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0C_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0C_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0C_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0C_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0C_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0C_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0C_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0C_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0C_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0C_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0C_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0C_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0C_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0C_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0C_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0C_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0C_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0C_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0C_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0C_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0C_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0C_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0C_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0C_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0D_Y0C_clk_out;
wire Tile_X0D_Y0C_clk_pass_through_out_bot;
wire Tile_X0D_Y0C_clk_pass_through_out_right;
wire [31:0] Tile_X0D_Y0C_config_out_config_addr;
wire [31:0] Tile_X0D_Y0C_config_out_config_data;
wire [0:0] Tile_X0D_Y0C_config_out_read;
wire [0:0] Tile_X0D_Y0C_config_out_write;
wire [8:0] Tile_X0D_Y0C_hi_unq1;
wire [7:0] Tile_X0D_Y0C_lo_unq1;
wire [31:0] Tile_X0D_Y0C_read_config_data;
wire Tile_X0D_Y0C_reset_out;
wire [0:0] Tile_X0D_Y0C_stall_out;
wire [8:0] Tile_X0D_Y0C_hi_out;
wire [7:0] Tile_X0D_Y0C_lo_out;
wire [15:0] Tile_X0D_Y0C_tile_id_in;
wire [0:0] Tile_X0D_Y0D_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0D_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0D_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0D_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0D_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0D_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0D_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0D_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0D_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0D_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0D_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0D_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0D_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0D_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0D_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0D_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0D_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0D_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0D_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0D_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0D_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0D_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0D_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0D_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0D_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0D_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0D_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0D_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0D_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0D_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0D_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0D_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0D_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0D_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0D_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0D_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0D_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0D_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0D_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0D_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0D_Y0D_clk_out;
wire Tile_X0D_Y0D_clk_pass_through_out_bot;
wire Tile_X0D_Y0D_clk_pass_through_out_right;
wire [31:0] Tile_X0D_Y0D_config_out_config_addr;
wire [31:0] Tile_X0D_Y0D_config_out_config_data;
wire [0:0] Tile_X0D_Y0D_config_out_read;
wire [0:0] Tile_X0D_Y0D_config_out_write;
wire [8:0] Tile_X0D_Y0D_hi_unq1;
wire [7:0] Tile_X0D_Y0D_lo_unq1;
wire [31:0] Tile_X0D_Y0D_read_config_data;
wire Tile_X0D_Y0D_reset_out;
wire [0:0] Tile_X0D_Y0D_stall_out;
wire [8:0] Tile_X0D_Y0D_hi_out;
wire [7:0] Tile_X0D_Y0D_lo_out;
wire [15:0] Tile_X0D_Y0D_tile_id_in;
wire [0:0] Tile_X0D_Y0E_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0E_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0E_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0E_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0E_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0E_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0E_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0E_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0E_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0E_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0E_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0E_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0E_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0E_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0E_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0E_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0E_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0E_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0E_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0E_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0E_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0E_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0E_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0E_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0E_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0E_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0E_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0E_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0E_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0E_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0E_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0E_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0E_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0E_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0E_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0E_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0E_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0E_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0E_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0E_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0D_Y0E_clk_out;
wire Tile_X0D_Y0E_clk_pass_through_out_bot;
wire Tile_X0D_Y0E_clk_pass_through_out_right;
wire [31:0] Tile_X0D_Y0E_config_out_config_addr;
wire [31:0] Tile_X0D_Y0E_config_out_config_data;
wire [0:0] Tile_X0D_Y0E_config_out_read;
wire [0:0] Tile_X0D_Y0E_config_out_write;
wire [8:0] Tile_X0D_Y0E_hi_unq1;
wire [7:0] Tile_X0D_Y0E_lo_unq1;
wire [31:0] Tile_X0D_Y0E_read_config_data;
wire Tile_X0D_Y0E_reset_out;
wire [0:0] Tile_X0D_Y0E_stall_out;
wire [8:0] Tile_X0D_Y0E_hi_out;
wire [7:0] Tile_X0D_Y0E_lo_out;
wire [15:0] Tile_X0D_Y0E_tile_id_in;
wire [0:0] Tile_X0D_Y0F_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0F_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0F_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0F_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0F_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0F_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0F_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0F_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0F_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0F_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0F_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0F_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0F_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0F_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0F_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0F_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0F_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0F_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0F_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0F_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0F_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0F_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0F_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0F_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0F_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0F_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0F_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0F_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0F_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0F_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0F_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0F_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0F_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0F_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0F_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0F_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0F_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0F_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y0F_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y0F_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0D_Y0F_clk_out;
wire Tile_X0D_Y0F_clk_pass_through_out_bot;
wire Tile_X0D_Y0F_clk_pass_through_out_right;
wire [31:0] Tile_X0D_Y0F_config_out_config_addr;
wire [31:0] Tile_X0D_Y0F_config_out_config_data;
wire [0:0] Tile_X0D_Y0F_config_out_read;
wire [0:0] Tile_X0D_Y0F_config_out_write;
wire [8:0] Tile_X0D_Y0F_hi_unq1;
wire [7:0] Tile_X0D_Y0F_lo_unq1;
wire [31:0] Tile_X0D_Y0F_read_config_data;
wire Tile_X0D_Y0F_reset_out;
wire [0:0] Tile_X0D_Y0F_stall_out;
wire [8:0] Tile_X0D_Y0F_hi_out;
wire [7:0] Tile_X0D_Y0F_lo_out;
wire [15:0] Tile_X0D_Y0F_tile_id_in;
wire [0:0] Tile_X0D_Y10_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y10_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y10_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y10_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y10_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y10_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y10_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y10_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y10_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y10_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y10_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y10_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y10_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y10_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y10_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y10_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y10_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y10_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y10_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y10_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y10_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y10_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y10_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y10_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y10_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y10_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y10_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y10_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y10_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y10_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y10_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y10_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y10_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y10_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0D_Y10_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y10_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y10_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0D_Y10_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0D_Y10_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0D_Y10_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0D_Y10_clk_out;
wire Tile_X0D_Y10_clk_pass_through_out_bot;
wire Tile_X0D_Y10_clk_pass_through_out_right;
wire [31:0] Tile_X0D_Y10_config_out_config_addr;
wire [31:0] Tile_X0D_Y10_config_out_config_data;
wire [0:0] Tile_X0D_Y10_config_out_read;
wire [0:0] Tile_X0D_Y10_config_out_write;
wire [8:0] Tile_X0D_Y10_hi_unq1;
wire [7:0] Tile_X0D_Y10_lo_unq1;
wire [31:0] Tile_X0D_Y10_read_config_data;
wire Tile_X0D_Y10_reset_out;
wire [0:0] Tile_X0D_Y10_stall_out;
wire [8:0] Tile_X0D_Y10_hi_out;
wire [7:0] Tile_X0D_Y10_lo_out;
wire [15:0] Tile_X0D_Y10_tile_id_in;
wire [0:0] Tile_X0E_Y00_io2glb_1;
wire [0:0] Tile_X0E_Y00_io2f_1;
wire [15:0] Tile_X0E_Y00_io2glb_16;
wire [15:0] Tile_X0E_Y00_io2f_16;
wire [8:0] Tile_X0E_Y00_hi;
wire [7:0] Tile_X0E_Y00_lo;
wire [0:0] Tile_X0E_Y01_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y01_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y01_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y01_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y01_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y01_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y01_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y01_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y01_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y01_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y01_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y01_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y01_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y01_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y01_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y01_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y01_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y01_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y01_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y01_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y01_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y01_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y01_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y01_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y01_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y01_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y01_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y01_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y01_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y01_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y01_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y01_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y01_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y01_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y01_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y01_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y01_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y01_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y01_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y01_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0E_Y01_clk_out;
wire Tile_X0E_Y01_clk_pass_through_out_bot;
wire Tile_X0E_Y01_clk_pass_through_out_right;
wire [31:0] Tile_X0E_Y01_config_out_config_addr;
wire [31:0] Tile_X0E_Y01_config_out_config_data;
wire [0:0] Tile_X0E_Y01_config_out_read;
wire [0:0] Tile_X0E_Y01_config_out_write;
wire [8:0] Tile_X0E_Y01_hi_unq1;
wire [7:0] Tile_X0E_Y01_lo_unq1;
wire [31:0] Tile_X0E_Y01_read_config_data;
wire Tile_X0E_Y01_reset_out;
wire [0:0] Tile_X0E_Y01_stall_out;
wire [8:0] Tile_X0E_Y01_hi_out;
wire [7:0] Tile_X0E_Y01_lo_out;
wire [15:0] Tile_X0E_Y01_tile_id_in;
wire [0:0] Tile_X0E_Y02_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y02_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y02_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y02_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y02_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y02_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y02_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y02_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y02_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y02_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y02_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y02_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y02_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y02_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y02_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y02_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y02_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y02_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y02_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y02_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y02_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y02_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y02_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y02_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y02_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y02_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y02_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y02_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y02_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y02_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y02_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y02_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y02_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y02_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y02_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y02_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y02_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y02_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y02_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y02_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0E_Y02_clk_out;
wire Tile_X0E_Y02_clk_pass_through_out_bot;
wire Tile_X0E_Y02_clk_pass_through_out_right;
wire [31:0] Tile_X0E_Y02_config_out_config_addr;
wire [31:0] Tile_X0E_Y02_config_out_config_data;
wire [0:0] Tile_X0E_Y02_config_out_read;
wire [0:0] Tile_X0E_Y02_config_out_write;
wire [8:0] Tile_X0E_Y02_hi_unq1;
wire [7:0] Tile_X0E_Y02_lo_unq1;
wire [31:0] Tile_X0E_Y02_read_config_data;
wire Tile_X0E_Y02_reset_out;
wire [0:0] Tile_X0E_Y02_stall_out;
wire [8:0] Tile_X0E_Y02_hi_out;
wire [7:0] Tile_X0E_Y02_lo_out;
wire [15:0] Tile_X0E_Y02_tile_id_in;
wire [0:0] Tile_X0E_Y03_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y03_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y03_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y03_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y03_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y03_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y03_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y03_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y03_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y03_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y03_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y03_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y03_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y03_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y03_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y03_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y03_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y03_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y03_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y03_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y03_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y03_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y03_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y03_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y03_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y03_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y03_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y03_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y03_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y03_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y03_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y03_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y03_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y03_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y03_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y03_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y03_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y03_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y03_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y03_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0E_Y03_clk_out;
wire Tile_X0E_Y03_clk_pass_through_out_bot;
wire Tile_X0E_Y03_clk_pass_through_out_right;
wire [31:0] Tile_X0E_Y03_config_out_config_addr;
wire [31:0] Tile_X0E_Y03_config_out_config_data;
wire [0:0] Tile_X0E_Y03_config_out_read;
wire [0:0] Tile_X0E_Y03_config_out_write;
wire [8:0] Tile_X0E_Y03_hi_unq1;
wire [7:0] Tile_X0E_Y03_lo_unq1;
wire [31:0] Tile_X0E_Y03_read_config_data;
wire Tile_X0E_Y03_reset_out;
wire [0:0] Tile_X0E_Y03_stall_out;
wire [8:0] Tile_X0E_Y03_hi_out;
wire [7:0] Tile_X0E_Y03_lo_out;
wire [15:0] Tile_X0E_Y03_tile_id_in;
wire [0:0] Tile_X0E_Y04_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y04_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y04_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y04_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y04_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y04_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y04_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y04_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y04_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y04_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y04_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y04_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y04_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y04_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y04_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y04_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y04_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y04_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y04_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y04_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y04_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y04_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y04_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y04_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y04_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y04_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y04_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y04_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y04_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y04_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y04_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y04_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y04_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y04_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y04_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y04_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y04_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y04_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y04_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y04_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0E_Y04_clk_out;
wire Tile_X0E_Y04_clk_pass_through_out_bot;
wire Tile_X0E_Y04_clk_pass_through_out_right;
wire [31:0] Tile_X0E_Y04_config_out_config_addr;
wire [31:0] Tile_X0E_Y04_config_out_config_data;
wire [0:0] Tile_X0E_Y04_config_out_read;
wire [0:0] Tile_X0E_Y04_config_out_write;
wire [8:0] Tile_X0E_Y04_hi_unq1;
wire [7:0] Tile_X0E_Y04_lo_unq1;
wire [31:0] Tile_X0E_Y04_read_config_data;
wire Tile_X0E_Y04_reset_out;
wire [0:0] Tile_X0E_Y04_stall_out;
wire [8:0] Tile_X0E_Y04_hi_out;
wire [7:0] Tile_X0E_Y04_lo_out;
wire [15:0] Tile_X0E_Y04_tile_id_in;
wire [0:0] Tile_X0E_Y05_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y05_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y05_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y05_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y05_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y05_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y05_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y05_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y05_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y05_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y05_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y05_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y05_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y05_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y05_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y05_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y05_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y05_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y05_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y05_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y05_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y05_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y05_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y05_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y05_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y05_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y05_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y05_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y05_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y05_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y05_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y05_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y05_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y05_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y05_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y05_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y05_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y05_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y05_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y05_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0E_Y05_clk_out;
wire Tile_X0E_Y05_clk_pass_through_out_bot;
wire Tile_X0E_Y05_clk_pass_through_out_right;
wire [31:0] Tile_X0E_Y05_config_out_config_addr;
wire [31:0] Tile_X0E_Y05_config_out_config_data;
wire [0:0] Tile_X0E_Y05_config_out_read;
wire [0:0] Tile_X0E_Y05_config_out_write;
wire [8:0] Tile_X0E_Y05_hi_unq1;
wire [7:0] Tile_X0E_Y05_lo_unq1;
wire [31:0] Tile_X0E_Y05_read_config_data;
wire Tile_X0E_Y05_reset_out;
wire [0:0] Tile_X0E_Y05_stall_out;
wire [8:0] Tile_X0E_Y05_hi_out;
wire [7:0] Tile_X0E_Y05_lo_out;
wire [15:0] Tile_X0E_Y05_tile_id_in;
wire [0:0] Tile_X0E_Y06_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y06_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y06_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y06_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y06_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y06_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y06_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y06_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y06_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y06_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y06_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y06_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y06_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y06_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y06_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y06_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y06_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y06_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y06_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y06_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y06_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y06_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y06_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y06_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y06_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y06_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y06_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y06_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y06_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y06_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y06_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y06_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y06_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y06_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y06_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y06_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y06_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y06_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y06_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y06_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0E_Y06_clk_out;
wire Tile_X0E_Y06_clk_pass_through_out_bot;
wire Tile_X0E_Y06_clk_pass_through_out_right;
wire [31:0] Tile_X0E_Y06_config_out_config_addr;
wire [31:0] Tile_X0E_Y06_config_out_config_data;
wire [0:0] Tile_X0E_Y06_config_out_read;
wire [0:0] Tile_X0E_Y06_config_out_write;
wire [8:0] Tile_X0E_Y06_hi_unq1;
wire [7:0] Tile_X0E_Y06_lo_unq1;
wire [31:0] Tile_X0E_Y06_read_config_data;
wire Tile_X0E_Y06_reset_out;
wire [0:0] Tile_X0E_Y06_stall_out;
wire [8:0] Tile_X0E_Y06_hi_out;
wire [7:0] Tile_X0E_Y06_lo_out;
wire [15:0] Tile_X0E_Y06_tile_id_in;
wire [0:0] Tile_X0E_Y07_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y07_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y07_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y07_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y07_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y07_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y07_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y07_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y07_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y07_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y07_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y07_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y07_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y07_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y07_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y07_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y07_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y07_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y07_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y07_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y07_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y07_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y07_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y07_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y07_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y07_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y07_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y07_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y07_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y07_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y07_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y07_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y07_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y07_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y07_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y07_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y07_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y07_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y07_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y07_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0E_Y07_clk_out;
wire Tile_X0E_Y07_clk_pass_through_out_bot;
wire Tile_X0E_Y07_clk_pass_through_out_right;
wire [31:0] Tile_X0E_Y07_config_out_config_addr;
wire [31:0] Tile_X0E_Y07_config_out_config_data;
wire [0:0] Tile_X0E_Y07_config_out_read;
wire [0:0] Tile_X0E_Y07_config_out_write;
wire [8:0] Tile_X0E_Y07_hi_unq1;
wire [7:0] Tile_X0E_Y07_lo_unq1;
wire [31:0] Tile_X0E_Y07_read_config_data;
wire Tile_X0E_Y07_reset_out;
wire [0:0] Tile_X0E_Y07_stall_out;
wire [8:0] Tile_X0E_Y07_hi_out;
wire [7:0] Tile_X0E_Y07_lo_out;
wire [15:0] Tile_X0E_Y07_tile_id_in;
wire [0:0] Tile_X0E_Y08_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y08_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y08_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y08_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y08_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y08_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y08_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y08_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y08_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y08_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y08_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y08_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y08_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y08_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y08_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y08_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y08_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y08_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y08_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y08_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y08_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y08_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y08_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y08_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y08_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y08_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y08_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y08_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y08_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y08_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y08_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y08_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y08_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y08_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y08_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y08_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y08_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y08_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y08_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y08_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0E_Y08_clk_out;
wire Tile_X0E_Y08_clk_pass_through_out_bot;
wire Tile_X0E_Y08_clk_pass_through_out_right;
wire [31:0] Tile_X0E_Y08_config_out_config_addr;
wire [31:0] Tile_X0E_Y08_config_out_config_data;
wire [0:0] Tile_X0E_Y08_config_out_read;
wire [0:0] Tile_X0E_Y08_config_out_write;
wire [8:0] Tile_X0E_Y08_hi_unq1;
wire [7:0] Tile_X0E_Y08_lo_unq1;
wire [31:0] Tile_X0E_Y08_read_config_data;
wire Tile_X0E_Y08_reset_out;
wire [0:0] Tile_X0E_Y08_stall_out;
wire [8:0] Tile_X0E_Y08_hi_out;
wire [7:0] Tile_X0E_Y08_lo_out;
wire [15:0] Tile_X0E_Y08_tile_id_in;
wire [0:0] Tile_X0E_Y09_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y09_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y09_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y09_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y09_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y09_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y09_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y09_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y09_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y09_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y09_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y09_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y09_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y09_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y09_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y09_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y09_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y09_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y09_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y09_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y09_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y09_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y09_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y09_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y09_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y09_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y09_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y09_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y09_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y09_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y09_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y09_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y09_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y09_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y09_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y09_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y09_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y09_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y09_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y09_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0E_Y09_clk_out;
wire Tile_X0E_Y09_clk_pass_through_out_bot;
wire Tile_X0E_Y09_clk_pass_through_out_right;
wire [31:0] Tile_X0E_Y09_config_out_config_addr;
wire [31:0] Tile_X0E_Y09_config_out_config_data;
wire [0:0] Tile_X0E_Y09_config_out_read;
wire [0:0] Tile_X0E_Y09_config_out_write;
wire [8:0] Tile_X0E_Y09_hi_unq1;
wire [7:0] Tile_X0E_Y09_lo_unq1;
wire [31:0] Tile_X0E_Y09_read_config_data;
wire Tile_X0E_Y09_reset_out;
wire [0:0] Tile_X0E_Y09_stall_out;
wire [8:0] Tile_X0E_Y09_hi_out;
wire [7:0] Tile_X0E_Y09_lo_out;
wire [15:0] Tile_X0E_Y09_tile_id_in;
wire [0:0] Tile_X0E_Y0A_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0A_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0A_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0A_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0A_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0A_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0A_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0A_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0A_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0A_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0A_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0A_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0A_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0A_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0A_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0A_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0A_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0A_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0A_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0A_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0A_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0A_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0A_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0A_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0A_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0A_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0A_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0A_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0A_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0A_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0A_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0A_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0A_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0A_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0A_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0A_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0A_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0A_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0A_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0A_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0E_Y0A_clk_out;
wire Tile_X0E_Y0A_clk_pass_through_out_bot;
wire Tile_X0E_Y0A_clk_pass_through_out_right;
wire [31:0] Tile_X0E_Y0A_config_out_config_addr;
wire [31:0] Tile_X0E_Y0A_config_out_config_data;
wire [0:0] Tile_X0E_Y0A_config_out_read;
wire [0:0] Tile_X0E_Y0A_config_out_write;
wire [8:0] Tile_X0E_Y0A_hi_unq1;
wire [7:0] Tile_X0E_Y0A_lo_unq1;
wire [31:0] Tile_X0E_Y0A_read_config_data;
wire Tile_X0E_Y0A_reset_out;
wire [0:0] Tile_X0E_Y0A_stall_out;
wire [8:0] Tile_X0E_Y0A_hi_out;
wire [7:0] Tile_X0E_Y0A_lo_out;
wire [15:0] Tile_X0E_Y0A_tile_id_in;
wire [0:0] Tile_X0E_Y0B_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0B_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0B_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0B_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0B_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0B_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0B_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0B_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0B_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0B_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0B_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0B_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0B_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0B_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0B_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0B_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0B_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0B_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0B_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0B_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0B_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0B_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0B_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0B_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0B_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0B_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0B_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0B_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0B_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0B_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0B_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0B_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0B_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0B_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0B_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0B_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0B_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0B_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0B_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0B_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0E_Y0B_clk_out;
wire Tile_X0E_Y0B_clk_pass_through_out_bot;
wire Tile_X0E_Y0B_clk_pass_through_out_right;
wire [31:0] Tile_X0E_Y0B_config_out_config_addr;
wire [31:0] Tile_X0E_Y0B_config_out_config_data;
wire [0:0] Tile_X0E_Y0B_config_out_read;
wire [0:0] Tile_X0E_Y0B_config_out_write;
wire [8:0] Tile_X0E_Y0B_hi_unq1;
wire [7:0] Tile_X0E_Y0B_lo_unq1;
wire [31:0] Tile_X0E_Y0B_read_config_data;
wire Tile_X0E_Y0B_reset_out;
wire [0:0] Tile_X0E_Y0B_stall_out;
wire [8:0] Tile_X0E_Y0B_hi_out;
wire [7:0] Tile_X0E_Y0B_lo_out;
wire [15:0] Tile_X0E_Y0B_tile_id_in;
wire [0:0] Tile_X0E_Y0C_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0C_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0C_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0C_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0C_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0C_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0C_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0C_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0C_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0C_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0C_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0C_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0C_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0C_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0C_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0C_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0C_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0C_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0C_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0C_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0C_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0C_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0C_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0C_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0C_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0C_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0C_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0C_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0C_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0C_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0C_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0C_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0C_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0C_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0C_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0C_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0C_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0C_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0C_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0C_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0E_Y0C_clk_out;
wire Tile_X0E_Y0C_clk_pass_through_out_bot;
wire Tile_X0E_Y0C_clk_pass_through_out_right;
wire [31:0] Tile_X0E_Y0C_config_out_config_addr;
wire [31:0] Tile_X0E_Y0C_config_out_config_data;
wire [0:0] Tile_X0E_Y0C_config_out_read;
wire [0:0] Tile_X0E_Y0C_config_out_write;
wire [8:0] Tile_X0E_Y0C_hi_unq1;
wire [7:0] Tile_X0E_Y0C_lo_unq1;
wire [31:0] Tile_X0E_Y0C_read_config_data;
wire Tile_X0E_Y0C_reset_out;
wire [0:0] Tile_X0E_Y0C_stall_out;
wire [8:0] Tile_X0E_Y0C_hi_out;
wire [7:0] Tile_X0E_Y0C_lo_out;
wire [15:0] Tile_X0E_Y0C_tile_id_in;
wire [0:0] Tile_X0E_Y0D_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0D_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0D_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0D_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0D_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0D_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0D_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0D_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0D_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0D_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0D_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0D_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0D_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0D_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0D_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0D_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0D_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0D_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0D_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0D_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0D_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0D_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0D_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0D_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0D_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0D_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0D_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0D_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0D_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0D_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0D_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0D_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0D_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0D_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0D_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0D_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0D_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0D_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0D_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0D_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0E_Y0D_clk_out;
wire Tile_X0E_Y0D_clk_pass_through_out_bot;
wire Tile_X0E_Y0D_clk_pass_through_out_right;
wire [31:0] Tile_X0E_Y0D_config_out_config_addr;
wire [31:0] Tile_X0E_Y0D_config_out_config_data;
wire [0:0] Tile_X0E_Y0D_config_out_read;
wire [0:0] Tile_X0E_Y0D_config_out_write;
wire [8:0] Tile_X0E_Y0D_hi_unq1;
wire [7:0] Tile_X0E_Y0D_lo_unq1;
wire [31:0] Tile_X0E_Y0D_read_config_data;
wire Tile_X0E_Y0D_reset_out;
wire [0:0] Tile_X0E_Y0D_stall_out;
wire [8:0] Tile_X0E_Y0D_hi_out;
wire [7:0] Tile_X0E_Y0D_lo_out;
wire [15:0] Tile_X0E_Y0D_tile_id_in;
wire [0:0] Tile_X0E_Y0E_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0E_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0E_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0E_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0E_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0E_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0E_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0E_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0E_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0E_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0E_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0E_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0E_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0E_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0E_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0E_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0E_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0E_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0E_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0E_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0E_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0E_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0E_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0E_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0E_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0E_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0E_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0E_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0E_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0E_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0E_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0E_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0E_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0E_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0E_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0E_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0E_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0E_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0E_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0E_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0E_Y0E_clk_out;
wire Tile_X0E_Y0E_clk_pass_through_out_bot;
wire Tile_X0E_Y0E_clk_pass_through_out_right;
wire [31:0] Tile_X0E_Y0E_config_out_config_addr;
wire [31:0] Tile_X0E_Y0E_config_out_config_data;
wire [0:0] Tile_X0E_Y0E_config_out_read;
wire [0:0] Tile_X0E_Y0E_config_out_write;
wire [8:0] Tile_X0E_Y0E_hi_unq1;
wire [7:0] Tile_X0E_Y0E_lo_unq1;
wire [31:0] Tile_X0E_Y0E_read_config_data;
wire Tile_X0E_Y0E_reset_out;
wire [0:0] Tile_X0E_Y0E_stall_out;
wire [8:0] Tile_X0E_Y0E_hi_out;
wire [7:0] Tile_X0E_Y0E_lo_out;
wire [15:0] Tile_X0E_Y0E_tile_id_in;
wire [0:0] Tile_X0E_Y0F_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0F_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0F_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0F_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0F_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0F_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0F_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0F_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0F_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0F_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0F_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0F_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0F_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0F_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0F_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0F_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0F_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0F_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0F_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0F_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0F_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0F_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0F_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0F_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0F_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0F_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0F_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0F_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0F_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0F_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0F_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0F_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0F_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0F_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0F_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0F_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0F_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0F_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y0F_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y0F_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0E_Y0F_clk_out;
wire Tile_X0E_Y0F_clk_pass_through_out_bot;
wire Tile_X0E_Y0F_clk_pass_through_out_right;
wire [31:0] Tile_X0E_Y0F_config_out_config_addr;
wire [31:0] Tile_X0E_Y0F_config_out_config_data;
wire [0:0] Tile_X0E_Y0F_config_out_read;
wire [0:0] Tile_X0E_Y0F_config_out_write;
wire [8:0] Tile_X0E_Y0F_hi_unq1;
wire [7:0] Tile_X0E_Y0F_lo_unq1;
wire [31:0] Tile_X0E_Y0F_read_config_data;
wire Tile_X0E_Y0F_reset_out;
wire [0:0] Tile_X0E_Y0F_stall_out;
wire [8:0] Tile_X0E_Y0F_hi_out;
wire [7:0] Tile_X0E_Y0F_lo_out;
wire [15:0] Tile_X0E_Y0F_tile_id_in;
wire [0:0] Tile_X0E_Y10_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y10_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y10_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y10_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y10_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y10_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y10_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y10_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y10_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y10_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y10_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y10_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y10_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y10_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y10_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y10_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y10_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y10_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y10_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y10_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y10_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y10_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y10_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y10_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y10_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y10_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y10_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y10_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y10_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y10_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y10_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y10_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y10_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y10_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0E_Y10_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y10_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y10_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0E_Y10_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0E_Y10_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0E_Y10_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0E_Y10_clk_out;
wire Tile_X0E_Y10_clk_pass_through_out_bot;
wire Tile_X0E_Y10_clk_pass_through_out_right;
wire [31:0] Tile_X0E_Y10_config_out_config_addr;
wire [31:0] Tile_X0E_Y10_config_out_config_data;
wire [0:0] Tile_X0E_Y10_config_out_read;
wire [0:0] Tile_X0E_Y10_config_out_write;
wire [8:0] Tile_X0E_Y10_hi_unq1;
wire [7:0] Tile_X0E_Y10_lo_unq1;
wire [31:0] Tile_X0E_Y10_read_config_data;
wire Tile_X0E_Y10_reset_out;
wire [0:0] Tile_X0E_Y10_stall_out;
wire [8:0] Tile_X0E_Y10_hi_out;
wire [7:0] Tile_X0E_Y10_lo_out;
wire [15:0] Tile_X0E_Y10_tile_id_in;
wire [0:0] Tile_X0F_Y00_io2glb_1;
wire [0:0] Tile_X0F_Y00_io2f_1;
wire [15:0] Tile_X0F_Y00_io2glb_16;
wire [15:0] Tile_X0F_Y00_io2f_16;
wire [8:0] Tile_X0F_Y00_hi;
wire [7:0] Tile_X0F_Y00_lo;
wire [0:0] Tile_X0F_Y01_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y01_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y01_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y01_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y01_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y01_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y01_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y01_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y01_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y01_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y01_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y01_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y01_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y01_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y01_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y01_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y01_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y01_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y01_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y01_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y01_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y01_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y01_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y01_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y01_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y01_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y01_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y01_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y01_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y01_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y01_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y01_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y01_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y01_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y01_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y01_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y01_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y01_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y01_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y01_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0F_Y01_clk_out;
wire [31:0] Tile_X0F_Y01_config_out_config_addr;
wire [31:0] Tile_X0F_Y01_config_out_config_data;
wire [0:0] Tile_X0F_Y01_config_out_read;
wire [0:0] Tile_X0F_Y01_config_out_write;
wire [8:0] Tile_X0F_Y01_hi_unq1;
wire [7:0] Tile_X0F_Y01_lo_unq1;
wire [31:0] Tile_X0F_Y01_read_config_data;
wire Tile_X0F_Y01_reset_out;
wire [0:0] Tile_X0F_Y01_stall_out;
wire [8:0] Tile_X0F_Y01_hi_out;
wire [7:0] Tile_X0F_Y01_lo_out;
wire [15:0] Tile_X0F_Y01_tile_id_in;
wire [0:0] Tile_X0F_Y02_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y02_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y02_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y02_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y02_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y02_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y02_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y02_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y02_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y02_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y02_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y02_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y02_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y02_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y02_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y02_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y02_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y02_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y02_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y02_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y02_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y02_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y02_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y02_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y02_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y02_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y02_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y02_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y02_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y02_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y02_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y02_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y02_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y02_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y02_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y02_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y02_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y02_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y02_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y02_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0F_Y02_clk_out;
wire [31:0] Tile_X0F_Y02_config_out_config_addr;
wire [31:0] Tile_X0F_Y02_config_out_config_data;
wire [0:0] Tile_X0F_Y02_config_out_read;
wire [0:0] Tile_X0F_Y02_config_out_write;
wire [8:0] Tile_X0F_Y02_hi_unq1;
wire [7:0] Tile_X0F_Y02_lo_unq1;
wire [31:0] Tile_X0F_Y02_read_config_data;
wire Tile_X0F_Y02_reset_out;
wire [0:0] Tile_X0F_Y02_stall_out;
wire [8:0] Tile_X0F_Y02_hi_out;
wire [7:0] Tile_X0F_Y02_lo_out;
wire [15:0] Tile_X0F_Y02_tile_id_in;
wire [0:0] Tile_X0F_Y03_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y03_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y03_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y03_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y03_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y03_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y03_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y03_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y03_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y03_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y03_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y03_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y03_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y03_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y03_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y03_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y03_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y03_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y03_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y03_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y03_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y03_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y03_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y03_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y03_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y03_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y03_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y03_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y03_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y03_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y03_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y03_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y03_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y03_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y03_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y03_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y03_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y03_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y03_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y03_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0F_Y03_clk_out;
wire [31:0] Tile_X0F_Y03_config_out_config_addr;
wire [31:0] Tile_X0F_Y03_config_out_config_data;
wire [0:0] Tile_X0F_Y03_config_out_read;
wire [0:0] Tile_X0F_Y03_config_out_write;
wire [8:0] Tile_X0F_Y03_hi_unq1;
wire [7:0] Tile_X0F_Y03_lo_unq1;
wire [31:0] Tile_X0F_Y03_read_config_data;
wire Tile_X0F_Y03_reset_out;
wire [0:0] Tile_X0F_Y03_stall_out;
wire [8:0] Tile_X0F_Y03_hi_out;
wire [7:0] Tile_X0F_Y03_lo_out;
wire [15:0] Tile_X0F_Y03_tile_id_in;
wire [0:0] Tile_X0F_Y04_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y04_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y04_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y04_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y04_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y04_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y04_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y04_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y04_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y04_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y04_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y04_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y04_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y04_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y04_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y04_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y04_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y04_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y04_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y04_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y04_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y04_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y04_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y04_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y04_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y04_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y04_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y04_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y04_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y04_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y04_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y04_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y04_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y04_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y04_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y04_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y04_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y04_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y04_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y04_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0F_Y04_clk_out;
wire [31:0] Tile_X0F_Y04_config_out_config_addr;
wire [31:0] Tile_X0F_Y04_config_out_config_data;
wire [0:0] Tile_X0F_Y04_config_out_read;
wire [0:0] Tile_X0F_Y04_config_out_write;
wire [8:0] Tile_X0F_Y04_hi_unq1;
wire [7:0] Tile_X0F_Y04_lo_unq1;
wire [31:0] Tile_X0F_Y04_read_config_data;
wire Tile_X0F_Y04_reset_out;
wire [0:0] Tile_X0F_Y04_stall_out;
wire [8:0] Tile_X0F_Y04_hi_out;
wire [7:0] Tile_X0F_Y04_lo_out;
wire [15:0] Tile_X0F_Y04_tile_id_in;
wire [0:0] Tile_X0F_Y05_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y05_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y05_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y05_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y05_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y05_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y05_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y05_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y05_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y05_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y05_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y05_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y05_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y05_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y05_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y05_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y05_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y05_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y05_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y05_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y05_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y05_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y05_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y05_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y05_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y05_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y05_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y05_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y05_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y05_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y05_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y05_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y05_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y05_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y05_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y05_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y05_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y05_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y05_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y05_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0F_Y05_clk_out;
wire [31:0] Tile_X0F_Y05_config_out_config_addr;
wire [31:0] Tile_X0F_Y05_config_out_config_data;
wire [0:0] Tile_X0F_Y05_config_out_read;
wire [0:0] Tile_X0F_Y05_config_out_write;
wire [8:0] Tile_X0F_Y05_hi_unq1;
wire [7:0] Tile_X0F_Y05_lo_unq1;
wire [31:0] Tile_X0F_Y05_read_config_data;
wire Tile_X0F_Y05_reset_out;
wire [0:0] Tile_X0F_Y05_stall_out;
wire [8:0] Tile_X0F_Y05_hi_out;
wire [7:0] Tile_X0F_Y05_lo_out;
wire [15:0] Tile_X0F_Y05_tile_id_in;
wire [0:0] Tile_X0F_Y06_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y06_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y06_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y06_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y06_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y06_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y06_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y06_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y06_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y06_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y06_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y06_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y06_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y06_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y06_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y06_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y06_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y06_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y06_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y06_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y06_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y06_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y06_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y06_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y06_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y06_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y06_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y06_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y06_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y06_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y06_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y06_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y06_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y06_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y06_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y06_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y06_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y06_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y06_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y06_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0F_Y06_clk_out;
wire [31:0] Tile_X0F_Y06_config_out_config_addr;
wire [31:0] Tile_X0F_Y06_config_out_config_data;
wire [0:0] Tile_X0F_Y06_config_out_read;
wire [0:0] Tile_X0F_Y06_config_out_write;
wire [8:0] Tile_X0F_Y06_hi_unq1;
wire [7:0] Tile_X0F_Y06_lo_unq1;
wire [31:0] Tile_X0F_Y06_read_config_data;
wire Tile_X0F_Y06_reset_out;
wire [0:0] Tile_X0F_Y06_stall_out;
wire [8:0] Tile_X0F_Y06_hi_out;
wire [7:0] Tile_X0F_Y06_lo_out;
wire [15:0] Tile_X0F_Y06_tile_id_in;
wire [0:0] Tile_X0F_Y07_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y07_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y07_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y07_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y07_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y07_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y07_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y07_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y07_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y07_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y07_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y07_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y07_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y07_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y07_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y07_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y07_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y07_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y07_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y07_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y07_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y07_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y07_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y07_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y07_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y07_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y07_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y07_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y07_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y07_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y07_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y07_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y07_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y07_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y07_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y07_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y07_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y07_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y07_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y07_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0F_Y07_clk_out;
wire [31:0] Tile_X0F_Y07_config_out_config_addr;
wire [31:0] Tile_X0F_Y07_config_out_config_data;
wire [0:0] Tile_X0F_Y07_config_out_read;
wire [0:0] Tile_X0F_Y07_config_out_write;
wire [8:0] Tile_X0F_Y07_hi_unq1;
wire [7:0] Tile_X0F_Y07_lo_unq1;
wire [31:0] Tile_X0F_Y07_read_config_data;
wire Tile_X0F_Y07_reset_out;
wire [0:0] Tile_X0F_Y07_stall_out;
wire [8:0] Tile_X0F_Y07_hi_out;
wire [7:0] Tile_X0F_Y07_lo_out;
wire [15:0] Tile_X0F_Y07_tile_id_in;
wire [0:0] Tile_X0F_Y08_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y08_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y08_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y08_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y08_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y08_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y08_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y08_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y08_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y08_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y08_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y08_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y08_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y08_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y08_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y08_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y08_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y08_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y08_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y08_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y08_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y08_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y08_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y08_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y08_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y08_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y08_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y08_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y08_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y08_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y08_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y08_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y08_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y08_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y08_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y08_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y08_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y08_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y08_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y08_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0F_Y08_clk_out;
wire [31:0] Tile_X0F_Y08_config_out_config_addr;
wire [31:0] Tile_X0F_Y08_config_out_config_data;
wire [0:0] Tile_X0F_Y08_config_out_read;
wire [0:0] Tile_X0F_Y08_config_out_write;
wire [8:0] Tile_X0F_Y08_hi_unq1;
wire [7:0] Tile_X0F_Y08_lo_unq1;
wire [31:0] Tile_X0F_Y08_read_config_data;
wire Tile_X0F_Y08_reset_out;
wire [0:0] Tile_X0F_Y08_stall_out;
wire [8:0] Tile_X0F_Y08_hi_out;
wire [7:0] Tile_X0F_Y08_lo_out;
wire [15:0] Tile_X0F_Y08_tile_id_in;
wire [0:0] Tile_X0F_Y09_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y09_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y09_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y09_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y09_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y09_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y09_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y09_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y09_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y09_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y09_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y09_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y09_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y09_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y09_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y09_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y09_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y09_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y09_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y09_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y09_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y09_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y09_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y09_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y09_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y09_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y09_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y09_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y09_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y09_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y09_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y09_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y09_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y09_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y09_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y09_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y09_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y09_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y09_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y09_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0F_Y09_clk_out;
wire [31:0] Tile_X0F_Y09_config_out_config_addr;
wire [31:0] Tile_X0F_Y09_config_out_config_data;
wire [0:0] Tile_X0F_Y09_config_out_read;
wire [0:0] Tile_X0F_Y09_config_out_write;
wire [8:0] Tile_X0F_Y09_hi_unq1;
wire [7:0] Tile_X0F_Y09_lo_unq1;
wire [31:0] Tile_X0F_Y09_read_config_data;
wire Tile_X0F_Y09_reset_out;
wire [0:0] Tile_X0F_Y09_stall_out;
wire [8:0] Tile_X0F_Y09_hi_out;
wire [7:0] Tile_X0F_Y09_lo_out;
wire [15:0] Tile_X0F_Y09_tile_id_in;
wire [0:0] Tile_X0F_Y0A_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0A_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0A_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0A_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0A_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0A_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0A_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0A_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0A_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0A_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0A_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0A_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0A_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0A_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0A_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0A_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0A_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0A_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0A_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0A_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0A_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0A_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0A_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0A_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0A_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0A_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0A_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0A_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0A_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0A_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0A_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0A_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0A_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0A_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0A_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0A_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0A_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0A_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0A_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0A_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0F_Y0A_clk_out;
wire [31:0] Tile_X0F_Y0A_config_out_config_addr;
wire [31:0] Tile_X0F_Y0A_config_out_config_data;
wire [0:0] Tile_X0F_Y0A_config_out_read;
wire [0:0] Tile_X0F_Y0A_config_out_write;
wire [8:0] Tile_X0F_Y0A_hi_unq1;
wire [7:0] Tile_X0F_Y0A_lo_unq1;
wire [31:0] Tile_X0F_Y0A_read_config_data;
wire Tile_X0F_Y0A_reset_out;
wire [0:0] Tile_X0F_Y0A_stall_out;
wire [8:0] Tile_X0F_Y0A_hi_out;
wire [7:0] Tile_X0F_Y0A_lo_out;
wire [15:0] Tile_X0F_Y0A_tile_id_in;
wire [0:0] Tile_X0F_Y0B_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0B_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0B_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0B_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0B_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0B_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0B_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0B_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0B_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0B_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0B_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0B_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0B_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0B_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0B_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0B_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0B_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0B_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0B_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0B_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0B_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0B_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0B_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0B_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0B_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0B_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0B_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0B_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0B_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0B_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0B_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0B_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0B_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0B_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0B_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0B_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0B_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0B_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0B_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0B_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0F_Y0B_clk_out;
wire [31:0] Tile_X0F_Y0B_config_out_config_addr;
wire [31:0] Tile_X0F_Y0B_config_out_config_data;
wire [0:0] Tile_X0F_Y0B_config_out_read;
wire [0:0] Tile_X0F_Y0B_config_out_write;
wire [8:0] Tile_X0F_Y0B_hi_unq1;
wire [7:0] Tile_X0F_Y0B_lo_unq1;
wire [31:0] Tile_X0F_Y0B_read_config_data;
wire Tile_X0F_Y0B_reset_out;
wire [0:0] Tile_X0F_Y0B_stall_out;
wire [8:0] Tile_X0F_Y0B_hi_out;
wire [7:0] Tile_X0F_Y0B_lo_out;
wire [15:0] Tile_X0F_Y0B_tile_id_in;
wire [0:0] Tile_X0F_Y0C_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0C_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0C_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0C_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0C_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0C_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0C_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0C_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0C_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0C_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0C_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0C_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0C_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0C_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0C_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0C_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0C_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0C_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0C_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0C_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0C_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0C_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0C_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0C_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0C_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0C_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0C_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0C_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0C_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0C_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0C_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0C_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0C_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0C_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0C_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0C_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0C_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0C_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0C_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0C_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0F_Y0C_clk_out;
wire [31:0] Tile_X0F_Y0C_config_out_config_addr;
wire [31:0] Tile_X0F_Y0C_config_out_config_data;
wire [0:0] Tile_X0F_Y0C_config_out_read;
wire [0:0] Tile_X0F_Y0C_config_out_write;
wire [8:0] Tile_X0F_Y0C_hi_unq1;
wire [7:0] Tile_X0F_Y0C_lo_unq1;
wire [31:0] Tile_X0F_Y0C_read_config_data;
wire Tile_X0F_Y0C_reset_out;
wire [0:0] Tile_X0F_Y0C_stall_out;
wire [8:0] Tile_X0F_Y0C_hi_out;
wire [7:0] Tile_X0F_Y0C_lo_out;
wire [15:0] Tile_X0F_Y0C_tile_id_in;
wire [0:0] Tile_X0F_Y0D_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0D_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0D_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0D_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0D_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0D_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0D_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0D_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0D_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0D_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0D_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0D_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0D_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0D_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0D_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0D_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0D_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0D_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0D_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0D_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0D_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0D_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0D_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0D_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0D_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0D_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0D_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0D_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0D_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0D_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0D_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0D_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0D_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0D_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0D_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0D_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0D_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0D_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0D_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0D_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0F_Y0D_clk_out;
wire [31:0] Tile_X0F_Y0D_config_out_config_addr;
wire [31:0] Tile_X0F_Y0D_config_out_config_data;
wire [0:0] Tile_X0F_Y0D_config_out_read;
wire [0:0] Tile_X0F_Y0D_config_out_write;
wire [8:0] Tile_X0F_Y0D_hi_unq1;
wire [7:0] Tile_X0F_Y0D_lo_unq1;
wire [31:0] Tile_X0F_Y0D_read_config_data;
wire Tile_X0F_Y0D_reset_out;
wire [0:0] Tile_X0F_Y0D_stall_out;
wire [8:0] Tile_X0F_Y0D_hi_out;
wire [7:0] Tile_X0F_Y0D_lo_out;
wire [15:0] Tile_X0F_Y0D_tile_id_in;
wire [0:0] Tile_X0F_Y0E_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0E_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0E_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0E_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0E_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0E_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0E_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0E_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0E_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0E_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0E_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0E_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0E_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0E_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0E_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0E_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0E_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0E_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0E_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0E_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0E_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0E_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0E_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0E_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0E_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0E_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0E_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0E_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0E_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0E_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0E_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0E_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0E_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0E_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0E_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0E_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0E_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0E_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0E_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0E_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0F_Y0E_clk_out;
wire [31:0] Tile_X0F_Y0E_config_out_config_addr;
wire [31:0] Tile_X0F_Y0E_config_out_config_data;
wire [0:0] Tile_X0F_Y0E_config_out_read;
wire [0:0] Tile_X0F_Y0E_config_out_write;
wire [8:0] Tile_X0F_Y0E_hi_unq1;
wire [7:0] Tile_X0F_Y0E_lo_unq1;
wire [31:0] Tile_X0F_Y0E_read_config_data;
wire Tile_X0F_Y0E_reset_out;
wire [0:0] Tile_X0F_Y0E_stall_out;
wire [8:0] Tile_X0F_Y0E_hi_out;
wire [7:0] Tile_X0F_Y0E_lo_out;
wire [15:0] Tile_X0F_Y0E_tile_id_in;
wire [0:0] Tile_X0F_Y0F_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0F_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0F_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0F_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0F_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0F_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0F_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0F_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0F_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0F_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0F_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0F_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0F_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0F_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0F_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0F_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0F_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0F_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0F_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0F_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0F_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0F_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0F_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0F_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0F_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0F_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0F_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0F_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0F_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0F_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0F_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0F_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0F_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0F_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0F_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0F_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0F_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0F_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y0F_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y0F_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0F_Y0F_clk_out;
wire [31:0] Tile_X0F_Y0F_config_out_config_addr;
wire [31:0] Tile_X0F_Y0F_config_out_config_data;
wire [0:0] Tile_X0F_Y0F_config_out_read;
wire [0:0] Tile_X0F_Y0F_config_out_write;
wire [8:0] Tile_X0F_Y0F_hi_unq1;
wire [7:0] Tile_X0F_Y0F_lo_unq1;
wire [31:0] Tile_X0F_Y0F_read_config_data;
wire Tile_X0F_Y0F_reset_out;
wire [0:0] Tile_X0F_Y0F_stall_out;
wire [8:0] Tile_X0F_Y0F_hi_out;
wire [7:0] Tile_X0F_Y0F_lo_out;
wire [15:0] Tile_X0F_Y0F_tile_id_in;
wire [0:0] Tile_X0F_Y10_SB_T0_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y10_SB_T0_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y10_SB_T0_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y10_SB_T0_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y10_SB_T0_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y10_SB_T0_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y10_SB_T0_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y10_SB_T0_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y10_SB_T1_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y10_SB_T1_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y10_SB_T1_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y10_SB_T1_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y10_SB_T1_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y10_SB_T1_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y10_SB_T1_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y10_SB_T1_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y10_SB_T2_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y10_SB_T2_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y10_SB_T2_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y10_SB_T2_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y10_SB_T2_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y10_SB_T2_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y10_SB_T2_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y10_SB_T2_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y10_SB_T3_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y10_SB_T3_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y10_SB_T3_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y10_SB_T3_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y10_SB_T3_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y10_SB_T3_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y10_SB_T3_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y10_SB_T3_WEST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y10_SB_T4_EAST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y10_SB_T4_EAST_SB_OUT_B16;
wire [0:0] Tile_X0F_Y10_SB_T4_NORTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y10_SB_T4_NORTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y10_SB_T4_SOUTH_SB_OUT_B1;
wire [15:0] Tile_X0F_Y10_SB_T4_SOUTH_SB_OUT_B16;
wire [0:0] Tile_X0F_Y10_SB_T4_WEST_SB_OUT_B1;
wire [15:0] Tile_X0F_Y10_SB_T4_WEST_SB_OUT_B16;
wire Tile_X0F_Y10_clk_out;
wire [31:0] Tile_X0F_Y10_config_out_config_addr;
wire [31:0] Tile_X0F_Y10_config_out_config_data;
wire [0:0] Tile_X0F_Y10_config_out_read;
wire [0:0] Tile_X0F_Y10_config_out_write;
wire [8:0] Tile_X0F_Y10_hi_unq1;
wire [7:0] Tile_X0F_Y10_lo_unq1;
wire [31:0] Tile_X0F_Y10_read_config_data;
wire Tile_X0F_Y10_reset_out;
wire [0:0] Tile_X0F_Y10_stall_out;
wire [8:0] Tile_X0F_Y10_hi_out;
wire [7:0] Tile_X0F_Y10_lo_out;
wire [15:0] Tile_X0F_Y10_tile_id_in;
wire [0:0] const_0_1_out;
wire [15:0] const_0_16_out;
wire [31:0] const_0_32_out;
wire [31:0] read_config_data_or_final_O;
ConfigPipeStage ConfigPipeStage_inst0 (
    .clk(Tile_X00_Y08_clk_out),
    .config_config_addr(Tile_X00_Y08_config_out_config_addr),
    .config_config_data(Tile_X00_Y08_config_out_config_data),
    .config_out_config_addr(ConfigPipeStage_inst0_config_out_config_addr),
    .config_out_config_data(ConfigPipeStage_inst0_config_out_config_data),
    .config_out_read(ConfigPipeStage_inst0_config_out_read),
    .config_out_write(ConfigPipeStage_inst0_config_out_write),
    .config_read(Tile_X00_Y08_config_out_read),
    .config_write(Tile_X00_Y08_config_out_write)
);
ConfigPipeStage ConfigPipeStage_inst1 (
    .clk(Tile_X01_Y08_clk_out),
    .config_config_addr(Tile_X01_Y08_config_out_config_addr),
    .config_config_data(Tile_X01_Y08_config_out_config_data),
    .config_out_config_addr(ConfigPipeStage_inst1_config_out_config_addr),
    .config_out_config_data(ConfigPipeStage_inst1_config_out_config_data),
    .config_out_read(ConfigPipeStage_inst1_config_out_read),
    .config_out_write(ConfigPipeStage_inst1_config_out_write),
    .config_read(Tile_X01_Y08_config_out_read),
    .config_write(Tile_X01_Y08_config_out_write)
);
ConfigPipeStage ConfigPipeStage_inst10 (
    .clk(Tile_X0A_Y08_clk_out),
    .config_config_addr(Tile_X0A_Y08_config_out_config_addr),
    .config_config_data(Tile_X0A_Y08_config_out_config_data),
    .config_out_config_addr(ConfigPipeStage_inst10_config_out_config_addr),
    .config_out_config_data(ConfigPipeStage_inst10_config_out_config_data),
    .config_out_read(ConfigPipeStage_inst10_config_out_read),
    .config_out_write(ConfigPipeStage_inst10_config_out_write),
    .config_read(Tile_X0A_Y08_config_out_read),
    .config_write(Tile_X0A_Y08_config_out_write)
);
ConfigPipeStage ConfigPipeStage_inst11 (
    .clk(Tile_X0B_Y08_clk_out),
    .config_config_addr(Tile_X0B_Y08_config_out_config_addr),
    .config_config_data(Tile_X0B_Y08_config_out_config_data),
    .config_out_config_addr(ConfigPipeStage_inst11_config_out_config_addr),
    .config_out_config_data(ConfigPipeStage_inst11_config_out_config_data),
    .config_out_read(ConfigPipeStage_inst11_config_out_read),
    .config_out_write(ConfigPipeStage_inst11_config_out_write),
    .config_read(Tile_X0B_Y08_config_out_read),
    .config_write(Tile_X0B_Y08_config_out_write)
);
ConfigPipeStage ConfigPipeStage_inst12 (
    .clk(Tile_X0C_Y08_clk_out),
    .config_config_addr(Tile_X0C_Y08_config_out_config_addr),
    .config_config_data(Tile_X0C_Y08_config_out_config_data),
    .config_out_config_addr(ConfigPipeStage_inst12_config_out_config_addr),
    .config_out_config_data(ConfigPipeStage_inst12_config_out_config_data),
    .config_out_read(ConfigPipeStage_inst12_config_out_read),
    .config_out_write(ConfigPipeStage_inst12_config_out_write),
    .config_read(Tile_X0C_Y08_config_out_read),
    .config_write(Tile_X0C_Y08_config_out_write)
);
ConfigPipeStage ConfigPipeStage_inst13 (
    .clk(Tile_X0D_Y08_clk_out),
    .config_config_addr(Tile_X0D_Y08_config_out_config_addr),
    .config_config_data(Tile_X0D_Y08_config_out_config_data),
    .config_out_config_addr(ConfigPipeStage_inst13_config_out_config_addr),
    .config_out_config_data(ConfigPipeStage_inst13_config_out_config_data),
    .config_out_read(ConfigPipeStage_inst13_config_out_read),
    .config_out_write(ConfigPipeStage_inst13_config_out_write),
    .config_read(Tile_X0D_Y08_config_out_read),
    .config_write(Tile_X0D_Y08_config_out_write)
);
ConfigPipeStage ConfigPipeStage_inst14 (
    .clk(Tile_X0E_Y08_clk_out),
    .config_config_addr(Tile_X0E_Y08_config_out_config_addr),
    .config_config_data(Tile_X0E_Y08_config_out_config_data),
    .config_out_config_addr(ConfigPipeStage_inst14_config_out_config_addr),
    .config_out_config_data(ConfigPipeStage_inst14_config_out_config_data),
    .config_out_read(ConfigPipeStage_inst14_config_out_read),
    .config_out_write(ConfigPipeStage_inst14_config_out_write),
    .config_read(Tile_X0E_Y08_config_out_read),
    .config_write(Tile_X0E_Y08_config_out_write)
);
ConfigPipeStage ConfigPipeStage_inst15 (
    .clk(Tile_X0F_Y08_clk_out),
    .config_config_addr(Tile_X0F_Y08_config_out_config_addr),
    .config_config_data(Tile_X0F_Y08_config_out_config_data),
    .config_out_config_addr(ConfigPipeStage_inst15_config_out_config_addr),
    .config_out_config_data(ConfigPipeStage_inst15_config_out_config_data),
    .config_out_read(ConfigPipeStage_inst15_config_out_read),
    .config_out_write(ConfigPipeStage_inst15_config_out_write),
    .config_read(Tile_X0F_Y08_config_out_read),
    .config_write(Tile_X0F_Y08_config_out_write)
);
ConfigPipeStage ConfigPipeStage_inst2 (
    .clk(Tile_X02_Y08_clk_out),
    .config_config_addr(Tile_X02_Y08_config_out_config_addr),
    .config_config_data(Tile_X02_Y08_config_out_config_data),
    .config_out_config_addr(ConfigPipeStage_inst2_config_out_config_addr),
    .config_out_config_data(ConfigPipeStage_inst2_config_out_config_data),
    .config_out_read(ConfigPipeStage_inst2_config_out_read),
    .config_out_write(ConfigPipeStage_inst2_config_out_write),
    .config_read(Tile_X02_Y08_config_out_read),
    .config_write(Tile_X02_Y08_config_out_write)
);
ConfigPipeStage ConfigPipeStage_inst3 (
    .clk(Tile_X03_Y08_clk_out),
    .config_config_addr(Tile_X03_Y08_config_out_config_addr),
    .config_config_data(Tile_X03_Y08_config_out_config_data),
    .config_out_config_addr(ConfigPipeStage_inst3_config_out_config_addr),
    .config_out_config_data(ConfigPipeStage_inst3_config_out_config_data),
    .config_out_read(ConfigPipeStage_inst3_config_out_read),
    .config_out_write(ConfigPipeStage_inst3_config_out_write),
    .config_read(Tile_X03_Y08_config_out_read),
    .config_write(Tile_X03_Y08_config_out_write)
);
ConfigPipeStage ConfigPipeStage_inst4 (
    .clk(Tile_X04_Y08_clk_out),
    .config_config_addr(Tile_X04_Y08_config_out_config_addr),
    .config_config_data(Tile_X04_Y08_config_out_config_data),
    .config_out_config_addr(ConfigPipeStage_inst4_config_out_config_addr),
    .config_out_config_data(ConfigPipeStage_inst4_config_out_config_data),
    .config_out_read(ConfigPipeStage_inst4_config_out_read),
    .config_out_write(ConfigPipeStage_inst4_config_out_write),
    .config_read(Tile_X04_Y08_config_out_read),
    .config_write(Tile_X04_Y08_config_out_write)
);
ConfigPipeStage ConfigPipeStage_inst5 (
    .clk(Tile_X05_Y08_clk_out),
    .config_config_addr(Tile_X05_Y08_config_out_config_addr),
    .config_config_data(Tile_X05_Y08_config_out_config_data),
    .config_out_config_addr(ConfigPipeStage_inst5_config_out_config_addr),
    .config_out_config_data(ConfigPipeStage_inst5_config_out_config_data),
    .config_out_read(ConfigPipeStage_inst5_config_out_read),
    .config_out_write(ConfigPipeStage_inst5_config_out_write),
    .config_read(Tile_X05_Y08_config_out_read),
    .config_write(Tile_X05_Y08_config_out_write)
);
ConfigPipeStage ConfigPipeStage_inst6 (
    .clk(Tile_X06_Y08_clk_out),
    .config_config_addr(Tile_X06_Y08_config_out_config_addr),
    .config_config_data(Tile_X06_Y08_config_out_config_data),
    .config_out_config_addr(ConfigPipeStage_inst6_config_out_config_addr),
    .config_out_config_data(ConfigPipeStage_inst6_config_out_config_data),
    .config_out_read(ConfigPipeStage_inst6_config_out_read),
    .config_out_write(ConfigPipeStage_inst6_config_out_write),
    .config_read(Tile_X06_Y08_config_out_read),
    .config_write(Tile_X06_Y08_config_out_write)
);
ConfigPipeStage ConfigPipeStage_inst7 (
    .clk(Tile_X07_Y08_clk_out),
    .config_config_addr(Tile_X07_Y08_config_out_config_addr),
    .config_config_data(Tile_X07_Y08_config_out_config_data),
    .config_out_config_addr(ConfigPipeStage_inst7_config_out_config_addr),
    .config_out_config_data(ConfigPipeStage_inst7_config_out_config_data),
    .config_out_read(ConfigPipeStage_inst7_config_out_read),
    .config_out_write(ConfigPipeStage_inst7_config_out_write),
    .config_read(Tile_X07_Y08_config_out_read),
    .config_write(Tile_X07_Y08_config_out_write)
);
ConfigPipeStage ConfigPipeStage_inst8 (
    .clk(Tile_X08_Y08_clk_out),
    .config_config_addr(Tile_X08_Y08_config_out_config_addr),
    .config_config_data(Tile_X08_Y08_config_out_config_data),
    .config_out_config_addr(ConfigPipeStage_inst8_config_out_config_addr),
    .config_out_config_data(ConfigPipeStage_inst8_config_out_config_data),
    .config_out_read(ConfigPipeStage_inst8_config_out_read),
    .config_out_write(ConfigPipeStage_inst8_config_out_write),
    .config_read(Tile_X08_Y08_config_out_read),
    .config_write(Tile_X08_Y08_config_out_write)
);
ConfigPipeStage ConfigPipeStage_inst9 (
    .clk(Tile_X09_Y08_clk_out),
    .config_config_addr(Tile_X09_Y08_config_out_config_addr),
    .config_config_data(Tile_X09_Y08_config_out_config_data),
    .config_out_config_addr(ConfigPipeStage_inst9_config_out_config_addr),
    .config_out_config_data(ConfigPipeStage_inst9_config_out_config_data),
    .config_out_read(ConfigPipeStage_inst9_config_out_read),
    .config_out_write(ConfigPipeStage_inst9_config_out_write),
    .config_read(Tile_X09_Y08_config_out_read),
    .config_write(Tile_X09_Y08_config_out_write)
);
wire [15:0] Tile_X00_Y00_tile_id;
assign Tile_X00_Y00_tile_id = {Tile_X00_Y00_lo[7],Tile_X00_Y00_lo[7:6],Tile_X00_Y00_lo[6:5],Tile_X00_Y00_lo[5:4],Tile_X00_Y00_lo[4:3],Tile_X00_Y00_lo[3:2],Tile_X00_Y00_lo[2:1],Tile_X00_Y00_lo[1:0],Tile_X00_Y00_lo[0]};
Tile_io_core Tile_X00_Y00 (
    .tile_id(Tile_X00_Y00_tile_id),
    .glb2io_1(glb2io_1_X00_Y00),
    .f2io_1(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B1),
    .io2glb_1(Tile_X00_Y00_io2glb_1),
    .io2f_1(Tile_X00_Y00_io2f_1),
    .glb2io_16(glb2io_16_X00_Y00),
    .f2io_16(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B16),
    .io2glb_16(Tile_X00_Y00_io2glb_16),
    .io2f_16(Tile_X00_Y00_io2f_16),
    .hi(Tile_X00_Y00_hi),
    .lo(Tile_X00_Y00_lo)
);
Tile_PE Tile_X00_Y01 (
    .SB_T0_EAST_SB_IN_B1(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X00_Y00_io2f_1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X00_Y00_io2f_16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y01_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(const_0_1_out),
    .SB_T0_WEST_SB_IN_B16(const_0_16_out),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X00_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X00_Y00_io2f_1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X00_Y00_io2f_16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y01_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(const_0_1_out),
    .SB_T1_WEST_SB_IN_B16(const_0_16_out),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X00_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X00_Y00_io2f_1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X00_Y00_io2f_16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y01_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(const_0_1_out),
    .SB_T2_WEST_SB_IN_B16(const_0_16_out),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X00_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X01_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X01_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X00_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X00_Y00_io2f_1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X00_Y00_io2f_16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y01_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X00_Y01_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(const_0_1_out),
    .SB_T3_WEST_SB_IN_B16(const_0_16_out),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X00_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X01_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X01_Y01_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X00_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X00_Y00_io2f_1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X00_Y00_io2f_16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y01_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X00_Y01_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(const_0_1_out),
    .SB_T4_WEST_SB_IN_B16(const_0_16_out),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X00_Y01_SB_T4_WEST_SB_OUT_B16),
    .clk(clk),
    .clk_out(Tile_X00_Y01_clk_out),
    .clk_pass_through(clk),
    .clk_pass_through_out_bot(Tile_X00_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X00_Y01_clk_pass_through_out_right),
    .config_config_addr(config_0_config_addr),
    .config_config_data(config_0_config_data),
    .config_out_config_addr(Tile_X00_Y01_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y01_config_out_config_data),
    .config_out_read(Tile_X00_Y01_config_out_read),
    .config_out_write(Tile_X00_Y01_config_out_write),
    .config_read(config_0_read),
    .config_write(config_0_write),
    .hi(Tile_X00_Y01_hi),
    .lo(Tile_X00_Y01_lo_unq1),
    .read_config_data(Tile_X00_Y01_read_config_data),
    .read_config_data_in(const_0_32_out),
    .reset(reset),
    .reset_out(Tile_X00_Y01_reset_out),
    .stall(stall[0]),
    .stall_out(Tile_X00_Y01_stall_out),
    .tile_id(Tile_X00_Y01_tile_id_in)
);
mantle_wire__typeBit8 Tile_X00_Y01_lo (
    .in(Tile_X00_Y01_lo_unq1),
    .out(Tile_X00_Y01_lo_out)
);
wire [15:0] Tile_X00_Y01_tile_id_out;
assign Tile_X00_Y01_tile_id_out = {Tile_X00_Y01_lo_out[7],Tile_X00_Y01_lo_out[7:6],Tile_X00_Y01_lo_out[6:5],Tile_X00_Y01_lo_out[5:4],Tile_X00_Y01_lo_out[4:3],Tile_X00_Y01_lo_out[3:2],Tile_X00_Y01_lo_out[2:1],Tile_X00_Y01_lo_out[1:0],Tile_X00_Y01_hi[0]};
mantle_wire__typeBitIn16 Tile_X00_Y01_tile_id (
    .in(Tile_X00_Y01_tile_id_in),
    .out(Tile_X00_Y01_tile_id_out)
);
Tile_PE Tile_X00_Y02 (
    .SB_T0_EAST_SB_IN_B1(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X00_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(const_0_1_out),
    .SB_T0_WEST_SB_IN_B16(const_0_16_out),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X00_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X00_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(const_0_1_out),
    .SB_T1_WEST_SB_IN_B16(const_0_16_out),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X00_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X00_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(const_0_1_out),
    .SB_T2_WEST_SB_IN_B16(const_0_16_out),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X00_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X01_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X01_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X00_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X00_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X00_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(const_0_1_out),
    .SB_T3_WEST_SB_IN_B16(const_0_16_out),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X00_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X01_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X01_Y02_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X00_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X00_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X00_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(const_0_1_out),
    .SB_T4_WEST_SB_IN_B16(const_0_16_out),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X00_Y02_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X00_Y01_clk_out),
    .clk_out(Tile_X00_Y02_clk_out),
    .clk_pass_through(Tile_X00_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X00_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X00_Y02_clk_pass_through_out_right),
    .config_config_addr(Tile_X00_Y01_config_out_config_addr),
    .config_config_data(Tile_X00_Y01_config_out_config_data),
    .config_out_config_addr(Tile_X00_Y02_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y02_config_out_config_data),
    .config_out_read(Tile_X00_Y02_config_out_read),
    .config_out_write(Tile_X00_Y02_config_out_write),
    .config_read(Tile_X00_Y01_config_out_read),
    .config_write(Tile_X00_Y01_config_out_write),
    .hi(Tile_X00_Y02_hi),
    .lo(Tile_X00_Y02_lo_unq1),
    .read_config_data(Tile_X00_Y02_read_config_data),
    .read_config_data_in(Tile_X00_Y01_read_config_data),
    .reset(Tile_X00_Y01_reset_out),
    .reset_out(Tile_X00_Y02_reset_out),
    .stall(Tile_X00_Y01_stall_out),
    .stall_out(Tile_X00_Y02_stall_out),
    .tile_id(Tile_X00_Y02_tile_id_in)
);
mantle_wire__typeBit8 Tile_X00_Y02_lo (
    .in(Tile_X00_Y02_lo_unq1),
    .out(Tile_X00_Y02_lo_out)
);
wire [15:0] Tile_X00_Y02_tile_id_out;
assign Tile_X00_Y02_tile_id_out = {Tile_X00_Y02_lo_out[7],Tile_X00_Y02_lo_out[7:6],Tile_X00_Y02_lo_out[6:5],Tile_X00_Y02_lo_out[5:4],Tile_X00_Y02_lo_out[4:3],Tile_X00_Y02_lo_out[3:2],Tile_X00_Y02_lo_out[2:1],Tile_X00_Y02_lo_out[1],Tile_X00_Y02_hi[1],Tile_X00_Y02_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X00_Y02_tile_id (
    .in(Tile_X00_Y02_tile_id_in),
    .out(Tile_X00_Y02_tile_id_out)
);
Tile_PE Tile_X00_Y03 (
    .SB_T0_EAST_SB_IN_B1(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X00_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(const_0_1_out),
    .SB_T0_WEST_SB_IN_B16(const_0_16_out),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X00_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X00_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(const_0_1_out),
    .SB_T1_WEST_SB_IN_B16(const_0_16_out),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X00_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X00_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(const_0_1_out),
    .SB_T2_WEST_SB_IN_B16(const_0_16_out),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X00_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X01_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X01_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X00_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X00_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X00_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(const_0_1_out),
    .SB_T3_WEST_SB_IN_B16(const_0_16_out),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X00_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X01_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X01_Y03_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X00_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X00_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X00_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(const_0_1_out),
    .SB_T4_WEST_SB_IN_B16(const_0_16_out),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X00_Y03_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X00_Y02_clk_out),
    .clk_out(Tile_X00_Y03_clk_out),
    .clk_pass_through(Tile_X00_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X00_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X00_Y03_clk_pass_through_out_right),
    .config_config_addr(Tile_X00_Y02_config_out_config_addr),
    .config_config_data(Tile_X00_Y02_config_out_config_data),
    .config_out_config_addr(Tile_X00_Y03_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y03_config_out_config_data),
    .config_out_read(Tile_X00_Y03_config_out_read),
    .config_out_write(Tile_X00_Y03_config_out_write),
    .config_read(Tile_X00_Y02_config_out_read),
    .config_write(Tile_X00_Y02_config_out_write),
    .hi(Tile_X00_Y03_hi_unq1),
    .lo(Tile_X00_Y03_lo_unq1),
    .read_config_data(Tile_X00_Y03_read_config_data),
    .read_config_data_in(Tile_X00_Y02_read_config_data),
    .reset(Tile_X00_Y02_reset_out),
    .reset_out(Tile_X00_Y03_reset_out),
    .stall(Tile_X00_Y02_stall_out),
    .stall_out(Tile_X00_Y03_stall_out),
    .tile_id(Tile_X00_Y03_tile_id_in)
);
mantle_wire__typeBit9 Tile_X00_Y03_hi (
    .in(Tile_X00_Y03_hi_unq1),
    .out(Tile_X00_Y03_hi_out)
);
mantle_wire__typeBit8 Tile_X00_Y03_lo (
    .in(Tile_X00_Y03_lo_unq1),
    .out(Tile_X00_Y03_lo_out)
);
wire [15:0] Tile_X00_Y03_tile_id_out;
assign Tile_X00_Y03_tile_id_out = {Tile_X00_Y03_lo_out[7],Tile_X00_Y03_lo_out[7:6],Tile_X00_Y03_lo_out[6:5],Tile_X00_Y03_lo_out[5:4],Tile_X00_Y03_lo_out[4:3],Tile_X00_Y03_lo_out[3:2],Tile_X00_Y03_lo_out[2:1],Tile_X00_Y03_lo_out[1],Tile_X00_Y03_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X00_Y03_tile_id (
    .in(Tile_X00_Y03_tile_id_in),
    .out(Tile_X00_Y03_tile_id_out)
);
Tile_PE Tile_X00_Y04 (
    .SB_T0_EAST_SB_IN_B1(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X00_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(const_0_1_out),
    .SB_T0_WEST_SB_IN_B16(const_0_16_out),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X00_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X00_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(const_0_1_out),
    .SB_T1_WEST_SB_IN_B16(const_0_16_out),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X00_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X00_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(const_0_1_out),
    .SB_T2_WEST_SB_IN_B16(const_0_16_out),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X00_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X01_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X01_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X00_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X00_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X00_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X00_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X00_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(const_0_1_out),
    .SB_T3_WEST_SB_IN_B16(const_0_16_out),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X00_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X01_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X01_Y04_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X00_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X00_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X00_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X00_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X00_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(const_0_1_out),
    .SB_T4_WEST_SB_IN_B16(const_0_16_out),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X00_Y04_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X00_Y03_clk_out),
    .clk_out(Tile_X00_Y04_clk_out),
    .clk_pass_through(Tile_X00_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X00_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X00_Y04_clk_pass_through_out_right),
    .config_config_addr(Tile_X00_Y03_config_out_config_addr),
    .config_config_data(Tile_X00_Y03_config_out_config_data),
    .config_out_config_addr(Tile_X00_Y04_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y04_config_out_config_data),
    .config_out_read(Tile_X00_Y04_config_out_read),
    .config_out_write(Tile_X00_Y04_config_out_write),
    .config_read(Tile_X00_Y03_config_out_read),
    .config_write(Tile_X00_Y03_config_out_write),
    .hi(Tile_X00_Y04_hi),
    .lo(Tile_X00_Y04_lo_unq1),
    .read_config_data(Tile_X00_Y04_read_config_data),
    .read_config_data_in(Tile_X00_Y03_read_config_data),
    .reset(Tile_X00_Y03_reset_out),
    .reset_out(Tile_X00_Y04_reset_out),
    .stall(Tile_X00_Y03_stall_out),
    .stall_out(Tile_X00_Y04_stall_out),
    .tile_id(Tile_X00_Y04_tile_id_in)
);
mantle_wire__typeBit8 Tile_X00_Y04_lo (
    .in(Tile_X00_Y04_lo_unq1),
    .out(Tile_X00_Y04_lo_out)
);
wire [15:0] Tile_X00_Y04_tile_id_out;
assign Tile_X00_Y04_tile_id_out = {Tile_X00_Y04_lo_out[7],Tile_X00_Y04_lo_out[7:6],Tile_X00_Y04_lo_out[6:5],Tile_X00_Y04_lo_out[5:4],Tile_X00_Y04_lo_out[4:3],Tile_X00_Y04_lo_out[3:2],Tile_X00_Y04_lo_out[2:1],Tile_X00_Y04_hi[1],Tile_X00_Y04_lo_out[0],Tile_X00_Y04_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X00_Y04_tile_id (
    .in(Tile_X00_Y04_tile_id_in),
    .out(Tile_X00_Y04_tile_id_out)
);
Tile_PE Tile_X00_Y05 (
    .SB_T0_EAST_SB_IN_B1(Tile_X01_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X01_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X00_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X00_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(const_0_1_out),
    .SB_T0_WEST_SB_IN_B16(const_0_16_out),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X00_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X01_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X01_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X00_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X00_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(const_0_1_out),
    .SB_T1_WEST_SB_IN_B16(const_0_16_out),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X00_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X01_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X01_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X00_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X00_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(const_0_1_out),
    .SB_T2_WEST_SB_IN_B16(const_0_16_out),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X00_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X01_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X01_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X00_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X00_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X00_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X00_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X00_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X00_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(const_0_1_out),
    .SB_T3_WEST_SB_IN_B16(const_0_16_out),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X00_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X01_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X01_Y05_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X00_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X00_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X00_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X00_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X00_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X00_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(const_0_1_out),
    .SB_T4_WEST_SB_IN_B16(const_0_16_out),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X00_Y05_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X00_Y04_clk_out),
    .clk_out(Tile_X00_Y05_clk_out),
    .clk_pass_through(Tile_X00_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X00_Y05_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X00_Y05_clk_pass_through_out_right),
    .config_config_addr(Tile_X00_Y04_config_out_config_addr),
    .config_config_data(Tile_X00_Y04_config_out_config_data),
    .config_out_config_addr(Tile_X00_Y05_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y05_config_out_config_data),
    .config_out_read(Tile_X00_Y05_config_out_read),
    .config_out_write(Tile_X00_Y05_config_out_write),
    .config_read(Tile_X00_Y04_config_out_read),
    .config_write(Tile_X00_Y04_config_out_write),
    .hi(Tile_X00_Y05_hi),
    .lo(Tile_X00_Y05_lo_unq1),
    .read_config_data(Tile_X00_Y05_read_config_data),
    .read_config_data_in(Tile_X00_Y04_read_config_data),
    .reset(Tile_X00_Y04_reset_out),
    .reset_out(Tile_X00_Y05_reset_out),
    .stall(Tile_X00_Y04_stall_out),
    .stall_out(Tile_X00_Y05_stall_out),
    .tile_id(Tile_X00_Y05_tile_id_in)
);
mantle_wire__typeBit8 Tile_X00_Y05_lo (
    .in(Tile_X00_Y05_lo_unq1),
    .out(Tile_X00_Y05_lo_out)
);
wire [15:0] Tile_X00_Y05_tile_id_out;
assign Tile_X00_Y05_tile_id_out = {Tile_X00_Y05_lo_out[7],Tile_X00_Y05_lo_out[7:6],Tile_X00_Y05_lo_out[6:5],Tile_X00_Y05_lo_out[5:4],Tile_X00_Y05_lo_out[4:3],Tile_X00_Y05_lo_out[3:2],Tile_X00_Y05_lo_out[2:1],Tile_X00_Y05_hi[1],Tile_X00_Y05_lo_out[0],Tile_X00_Y05_hi[0]};
mantle_wire__typeBitIn16 Tile_X00_Y05_tile_id (
    .in(Tile_X00_Y05_tile_id_in),
    .out(Tile_X00_Y05_tile_id_out)
);
Tile_PE Tile_X00_Y06 (
    .SB_T0_EAST_SB_IN_B1(Tile_X01_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X01_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X00_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X00_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X00_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(const_0_1_out),
    .SB_T0_WEST_SB_IN_B16(const_0_16_out),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X00_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X01_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X01_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X00_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X00_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X00_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(const_0_1_out),
    .SB_T1_WEST_SB_IN_B16(const_0_16_out),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X00_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X01_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X01_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X00_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X00_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X00_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(const_0_1_out),
    .SB_T2_WEST_SB_IN_B16(const_0_16_out),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X00_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X01_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X01_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X00_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X00_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X00_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X00_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X00_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X00_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X00_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(const_0_1_out),
    .SB_T3_WEST_SB_IN_B16(const_0_16_out),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X00_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X01_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X01_Y06_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X00_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X00_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X00_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X00_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X00_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X00_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X00_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(const_0_1_out),
    .SB_T4_WEST_SB_IN_B16(const_0_16_out),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X00_Y06_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X00_Y05_clk_out),
    .clk_out(Tile_X00_Y06_clk_out),
    .clk_pass_through(Tile_X00_Y05_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X00_Y06_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X00_Y06_clk_pass_through_out_right),
    .config_config_addr(Tile_X00_Y05_config_out_config_addr),
    .config_config_data(Tile_X00_Y05_config_out_config_data),
    .config_out_config_addr(Tile_X00_Y06_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y06_config_out_config_data),
    .config_out_read(Tile_X00_Y06_config_out_read),
    .config_out_write(Tile_X00_Y06_config_out_write),
    .config_read(Tile_X00_Y05_config_out_read),
    .config_write(Tile_X00_Y05_config_out_write),
    .hi(Tile_X00_Y06_hi),
    .lo(Tile_X00_Y06_lo_unq1),
    .read_config_data(Tile_X00_Y06_read_config_data),
    .read_config_data_in(Tile_X00_Y05_read_config_data),
    .reset(Tile_X00_Y05_reset_out),
    .reset_out(Tile_X00_Y06_reset_out),
    .stall(Tile_X00_Y05_stall_out),
    .stall_out(Tile_X00_Y06_stall_out),
    .tile_id(Tile_X00_Y06_tile_id_in)
);
mantle_wire__typeBit8 Tile_X00_Y06_lo (
    .in(Tile_X00_Y06_lo_unq1),
    .out(Tile_X00_Y06_lo_out)
);
wire [15:0] Tile_X00_Y06_tile_id_out;
assign Tile_X00_Y06_tile_id_out = {Tile_X00_Y06_lo_out[7],Tile_X00_Y06_lo_out[7:6],Tile_X00_Y06_lo_out[6:5],Tile_X00_Y06_lo_out[5:4],Tile_X00_Y06_lo_out[4:3],Tile_X00_Y06_lo_out[3:2],Tile_X00_Y06_lo_out[2:1],Tile_X00_Y06_hi[1],Tile_X00_Y06_hi[1],Tile_X00_Y06_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X00_Y06_tile_id (
    .in(Tile_X00_Y06_tile_id_in),
    .out(Tile_X00_Y06_tile_id_out)
);
Tile_PE Tile_X00_Y07 (
    .SB_T0_EAST_SB_IN_B1(Tile_X01_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X01_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X00_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X00_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X00_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(const_0_1_out),
    .SB_T0_WEST_SB_IN_B16(const_0_16_out),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X00_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X01_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X01_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X00_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X00_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X00_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(const_0_1_out),
    .SB_T1_WEST_SB_IN_B16(const_0_16_out),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X00_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X01_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X01_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X00_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X00_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X00_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(const_0_1_out),
    .SB_T2_WEST_SB_IN_B16(const_0_16_out),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X00_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X01_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X01_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X00_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X00_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X00_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X00_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X00_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X00_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X00_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(const_0_1_out),
    .SB_T3_WEST_SB_IN_B16(const_0_16_out),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X00_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X01_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X01_Y07_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X00_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X00_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X00_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X00_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X00_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X00_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X00_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(const_0_1_out),
    .SB_T4_WEST_SB_IN_B16(const_0_16_out),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X00_Y07_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X00_Y06_clk_out),
    .clk_out(Tile_X00_Y07_clk_out),
    .clk_pass_through(Tile_X00_Y06_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X00_Y07_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X00_Y07_clk_pass_through_out_right),
    .config_config_addr(Tile_X00_Y06_config_out_config_addr),
    .config_config_data(Tile_X00_Y06_config_out_config_data),
    .config_out_config_addr(Tile_X00_Y07_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y07_config_out_config_data),
    .config_out_read(Tile_X00_Y07_config_out_read),
    .config_out_write(Tile_X00_Y07_config_out_write),
    .config_read(Tile_X00_Y06_config_out_read),
    .config_write(Tile_X00_Y06_config_out_write),
    .hi(Tile_X00_Y07_hi_unq1),
    .lo(Tile_X00_Y07_lo_unq1),
    .read_config_data(Tile_X00_Y07_read_config_data),
    .read_config_data_in(Tile_X00_Y06_read_config_data),
    .reset(Tile_X00_Y06_reset_out),
    .reset_out(Tile_X00_Y07_reset_out),
    .stall(Tile_X00_Y06_stall_out),
    .stall_out(Tile_X00_Y07_stall_out),
    .tile_id(Tile_X00_Y07_tile_id_in)
);
mantle_wire__typeBit9 Tile_X00_Y07_hi (
    .in(Tile_X00_Y07_hi_unq1),
    .out(Tile_X00_Y07_hi_out)
);
mantle_wire__typeBit8 Tile_X00_Y07_lo (
    .in(Tile_X00_Y07_lo_unq1),
    .out(Tile_X00_Y07_lo_out)
);
wire [15:0] Tile_X00_Y07_tile_id_out;
assign Tile_X00_Y07_tile_id_out = {Tile_X00_Y07_lo_out[7],Tile_X00_Y07_lo_out[7:6],Tile_X00_Y07_lo_out[6:5],Tile_X00_Y07_lo_out[5:4],Tile_X00_Y07_lo_out[4:3],Tile_X00_Y07_lo_out[3:2],Tile_X00_Y07_lo_out[2:1],Tile_X00_Y07_hi_out[1],Tile_X00_Y07_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X00_Y07_tile_id (
    .in(Tile_X00_Y07_tile_id_in),
    .out(Tile_X00_Y07_tile_id_out)
);
Tile_PE Tile_X00_Y08 (
    .SB_T0_EAST_SB_IN_B1(Tile_X01_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X01_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X00_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X00_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X00_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(const_0_1_out),
    .SB_T0_WEST_SB_IN_B16(const_0_16_out),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X00_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X01_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X01_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X00_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X00_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X00_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(const_0_1_out),
    .SB_T1_WEST_SB_IN_B16(const_0_16_out),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X00_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X01_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X01_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X00_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X00_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X00_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(const_0_1_out),
    .SB_T2_WEST_SB_IN_B16(const_0_16_out),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X00_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X01_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X01_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X00_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X00_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X00_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X00_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X00_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X00_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X00_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(const_0_1_out),
    .SB_T3_WEST_SB_IN_B16(const_0_16_out),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X00_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X01_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X01_Y08_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X00_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X00_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X00_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X00_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X00_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X00_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X00_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(const_0_1_out),
    .SB_T4_WEST_SB_IN_B16(const_0_16_out),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X00_Y08_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X00_Y07_clk_out),
    .clk_out(Tile_X00_Y08_clk_out),
    .clk_pass_through(Tile_X00_Y07_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X00_Y08_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X00_Y08_clk_pass_through_out_right),
    .config_config_addr(Tile_X00_Y07_config_out_config_addr),
    .config_config_data(Tile_X00_Y07_config_out_config_data),
    .config_out_config_addr(Tile_X00_Y08_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y08_config_out_config_data),
    .config_out_read(Tile_X00_Y08_config_out_read),
    .config_out_write(Tile_X00_Y08_config_out_write),
    .config_read(Tile_X00_Y07_config_out_read),
    .config_write(Tile_X00_Y07_config_out_write),
    .hi(Tile_X00_Y08_hi),
    .lo(Tile_X00_Y08_lo_unq1),
    .read_config_data(Tile_X00_Y08_read_config_data),
    .read_config_data_in(Tile_X00_Y07_read_config_data),
    .reset(Tile_X00_Y07_reset_out),
    .reset_out(Tile_X00_Y08_reset_out),
    .stall(Tile_X00_Y07_stall_out),
    .stall_out(Tile_X00_Y08_stall_out),
    .tile_id(Tile_X00_Y08_tile_id_in)
);
mantle_wire__typeBit8 Tile_X00_Y08_lo (
    .in(Tile_X00_Y08_lo_unq1),
    .out(Tile_X00_Y08_lo_out)
);
wire [15:0] Tile_X00_Y08_tile_id_out;
assign Tile_X00_Y08_tile_id_out = {Tile_X00_Y08_lo_out[7],Tile_X00_Y08_lo_out[7:6],Tile_X00_Y08_lo_out[6:5],Tile_X00_Y08_lo_out[5:4],Tile_X00_Y08_lo_out[4:3],Tile_X00_Y08_lo_out[3:2],Tile_X00_Y08_lo_out[2],Tile_X00_Y08_hi[2],Tile_X00_Y08_lo_out[1:0],Tile_X00_Y08_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X00_Y08_tile_id (
    .in(Tile_X00_Y08_tile_id_in),
    .out(Tile_X00_Y08_tile_id_out)
);
Tile_PE Tile_X00_Y09 (
    .SB_T0_EAST_SB_IN_B1(Tile_X01_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X01_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X00_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X00_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X00_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(const_0_1_out),
    .SB_T0_WEST_SB_IN_B16(const_0_16_out),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X00_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X01_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X01_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X00_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X00_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X00_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(const_0_1_out),
    .SB_T1_WEST_SB_IN_B16(const_0_16_out),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X00_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X01_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X01_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X00_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X00_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X00_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(const_0_1_out),
    .SB_T2_WEST_SB_IN_B16(const_0_16_out),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X00_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X01_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X01_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X00_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X00_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X00_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X00_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X00_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X00_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X00_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(const_0_1_out),
    .SB_T3_WEST_SB_IN_B16(const_0_16_out),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X00_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X01_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X01_Y09_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X00_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X00_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X00_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X00_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X00_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X00_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X00_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(const_0_1_out),
    .SB_T4_WEST_SB_IN_B16(const_0_16_out),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X00_Y09_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X00_Y08_clk_out),
    .clk_out(Tile_X00_Y09_clk_out),
    .clk_pass_through(Tile_X00_Y08_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X00_Y09_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X00_Y09_clk_pass_through_out_right),
    .config_config_addr(ConfigPipeStage_inst0_config_out_config_addr),
    .config_config_data(ConfigPipeStage_inst0_config_out_config_data),
    .config_out_config_addr(Tile_X00_Y09_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y09_config_out_config_data),
    .config_out_read(Tile_X00_Y09_config_out_read),
    .config_out_write(Tile_X00_Y09_config_out_write),
    .config_read(ConfigPipeStage_inst0_config_out_read),
    .config_write(ConfigPipeStage_inst0_config_out_write),
    .hi(Tile_X00_Y09_hi),
    .lo(Tile_X00_Y09_lo_unq1),
    .read_config_data(Tile_X00_Y09_read_config_data),
    .read_config_data_in(Tile_X00_Y08_read_config_data),
    .reset(Tile_X00_Y08_reset_out),
    .reset_out(Tile_X00_Y09_reset_out),
    .stall(Tile_X00_Y08_stall_out),
    .stall_out(Tile_X00_Y09_stall_out),
    .tile_id(Tile_X00_Y09_tile_id_in)
);
mantle_wire__typeBit8 Tile_X00_Y09_lo (
    .in(Tile_X00_Y09_lo_unq1),
    .out(Tile_X00_Y09_lo_out)
);
wire [15:0] Tile_X00_Y09_tile_id_out;
assign Tile_X00_Y09_tile_id_out = {Tile_X00_Y09_lo_out[7],Tile_X00_Y09_lo_out[7:6],Tile_X00_Y09_lo_out[6:5],Tile_X00_Y09_lo_out[5:4],Tile_X00_Y09_lo_out[4:3],Tile_X00_Y09_lo_out[3:2],Tile_X00_Y09_lo_out[2],Tile_X00_Y09_hi[2],Tile_X00_Y09_lo_out[1:0],Tile_X00_Y09_hi[0]};
mantle_wire__typeBitIn16 Tile_X00_Y09_tile_id (
    .in(Tile_X00_Y09_tile_id_in),
    .out(Tile_X00_Y09_tile_id_out)
);
Tile_PE Tile_X00_Y0A (
    .SB_T0_EAST_SB_IN_B1(Tile_X01_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X01_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X00_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X00_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X00_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(const_0_1_out),
    .SB_T0_WEST_SB_IN_B16(const_0_16_out),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X00_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X01_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X01_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X00_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X00_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X00_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(const_0_1_out),
    .SB_T1_WEST_SB_IN_B16(const_0_16_out),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X00_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X01_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X01_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X00_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X00_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X00_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(const_0_1_out),
    .SB_T2_WEST_SB_IN_B16(const_0_16_out),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X00_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X01_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X01_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X00_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X00_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X00_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X00_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X00_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X00_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X00_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(const_0_1_out),
    .SB_T3_WEST_SB_IN_B16(const_0_16_out),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X00_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X01_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X01_Y0A_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X00_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X00_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X00_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X00_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X00_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X00_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X00_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(const_0_1_out),
    .SB_T4_WEST_SB_IN_B16(const_0_16_out),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X00_Y0A_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X00_Y09_clk_out),
    .clk_out(Tile_X00_Y0A_clk_out),
    .clk_pass_through(Tile_X00_Y09_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X00_Y0A_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X00_Y0A_clk_pass_through_out_right),
    .config_config_addr(Tile_X00_Y09_config_out_config_addr),
    .config_config_data(Tile_X00_Y09_config_out_config_data),
    .config_out_config_addr(Tile_X00_Y0A_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y0A_config_out_config_data),
    .config_out_read(Tile_X00_Y0A_config_out_read),
    .config_out_write(Tile_X00_Y0A_config_out_write),
    .config_read(Tile_X00_Y09_config_out_read),
    .config_write(Tile_X00_Y09_config_out_write),
    .hi(Tile_X00_Y0A_hi),
    .lo(Tile_X00_Y0A_lo_unq1),
    .read_config_data(Tile_X00_Y0A_read_config_data),
    .read_config_data_in(Tile_X00_Y09_read_config_data),
    .reset(Tile_X00_Y09_reset_out),
    .reset_out(Tile_X00_Y0A_reset_out),
    .stall(Tile_X00_Y09_stall_out),
    .stall_out(Tile_X00_Y0A_stall_out),
    .tile_id(Tile_X00_Y0A_tile_id_in)
);
mantle_wire__typeBit8 Tile_X00_Y0A_lo (
    .in(Tile_X00_Y0A_lo_unq1),
    .out(Tile_X00_Y0A_lo_out)
);
wire [15:0] Tile_X00_Y0A_tile_id_out;
assign Tile_X00_Y0A_tile_id_out = {Tile_X00_Y0A_lo_out[7],Tile_X00_Y0A_lo_out[7:6],Tile_X00_Y0A_lo_out[6:5],Tile_X00_Y0A_lo_out[5:4],Tile_X00_Y0A_lo_out[4:3],Tile_X00_Y0A_lo_out[3:2],Tile_X00_Y0A_lo_out[2],Tile_X00_Y0A_hi[2],Tile_X00_Y0A_lo_out[1],Tile_X00_Y0A_hi[1],Tile_X00_Y0A_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X00_Y0A_tile_id (
    .in(Tile_X00_Y0A_tile_id_in),
    .out(Tile_X00_Y0A_tile_id_out)
);
Tile_PE Tile_X00_Y0B (
    .SB_T0_EAST_SB_IN_B1(Tile_X01_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X01_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X00_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X00_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X00_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(const_0_1_out),
    .SB_T0_WEST_SB_IN_B16(const_0_16_out),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X00_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X01_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X01_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X00_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X00_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X00_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(const_0_1_out),
    .SB_T1_WEST_SB_IN_B16(const_0_16_out),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X00_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X01_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X01_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X00_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X00_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X00_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(const_0_1_out),
    .SB_T2_WEST_SB_IN_B16(const_0_16_out),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X00_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X01_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X01_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X00_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X00_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X00_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X00_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X00_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X00_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X00_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(const_0_1_out),
    .SB_T3_WEST_SB_IN_B16(const_0_16_out),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X00_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X01_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X01_Y0B_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X00_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X00_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X00_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X00_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X00_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X00_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X00_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(const_0_1_out),
    .SB_T4_WEST_SB_IN_B16(const_0_16_out),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X00_Y0B_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X00_Y0A_clk_out),
    .clk_out(Tile_X00_Y0B_clk_out),
    .clk_pass_through(Tile_X00_Y0A_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X00_Y0B_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X00_Y0B_clk_pass_through_out_right),
    .config_config_addr(Tile_X00_Y0A_config_out_config_addr),
    .config_config_data(Tile_X00_Y0A_config_out_config_data),
    .config_out_config_addr(Tile_X00_Y0B_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y0B_config_out_config_data),
    .config_out_read(Tile_X00_Y0B_config_out_read),
    .config_out_write(Tile_X00_Y0B_config_out_write),
    .config_read(Tile_X00_Y0A_config_out_read),
    .config_write(Tile_X00_Y0A_config_out_write),
    .hi(Tile_X00_Y0B_hi_unq1),
    .lo(Tile_X00_Y0B_lo_unq1),
    .read_config_data(Tile_X00_Y0B_read_config_data),
    .read_config_data_in(Tile_X00_Y0A_read_config_data),
    .reset(Tile_X00_Y0A_reset_out),
    .reset_out(Tile_X00_Y0B_reset_out),
    .stall(Tile_X00_Y0A_stall_out),
    .stall_out(Tile_X00_Y0B_stall_out),
    .tile_id(Tile_X00_Y0B_tile_id_in)
);
mantle_wire__typeBit9 Tile_X00_Y0B_hi (
    .in(Tile_X00_Y0B_hi_unq1),
    .out(Tile_X00_Y0B_hi_out)
);
mantle_wire__typeBit8 Tile_X00_Y0B_lo (
    .in(Tile_X00_Y0B_lo_unq1),
    .out(Tile_X00_Y0B_lo_out)
);
wire [15:0] Tile_X00_Y0B_tile_id_out;
assign Tile_X00_Y0B_tile_id_out = {Tile_X00_Y0B_lo_out[7],Tile_X00_Y0B_lo_out[7:6],Tile_X00_Y0B_lo_out[6:5],Tile_X00_Y0B_lo_out[5:4],Tile_X00_Y0B_lo_out[4:3],Tile_X00_Y0B_lo_out[3:2],Tile_X00_Y0B_lo_out[2],Tile_X00_Y0B_hi_out[2],Tile_X00_Y0B_lo_out[1],Tile_X00_Y0B_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X00_Y0B_tile_id (
    .in(Tile_X00_Y0B_tile_id_in),
    .out(Tile_X00_Y0B_tile_id_out)
);
Tile_PE Tile_X00_Y0C (
    .SB_T0_EAST_SB_IN_B1(Tile_X01_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X01_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X00_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X00_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X00_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(const_0_1_out),
    .SB_T0_WEST_SB_IN_B16(const_0_16_out),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X00_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X01_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X01_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X00_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X00_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X00_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(const_0_1_out),
    .SB_T1_WEST_SB_IN_B16(const_0_16_out),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X00_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X01_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X01_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X00_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X00_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X00_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(const_0_1_out),
    .SB_T2_WEST_SB_IN_B16(const_0_16_out),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X00_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X01_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X01_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X00_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X00_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X00_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X00_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X00_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X00_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X00_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(const_0_1_out),
    .SB_T3_WEST_SB_IN_B16(const_0_16_out),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X00_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X01_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X01_Y0C_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X00_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X00_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X00_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X00_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X00_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X00_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X00_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(const_0_1_out),
    .SB_T4_WEST_SB_IN_B16(const_0_16_out),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X00_Y0C_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X00_Y0B_clk_out),
    .clk_out(Tile_X00_Y0C_clk_out),
    .clk_pass_through(Tile_X00_Y0B_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X00_Y0C_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X00_Y0C_clk_pass_through_out_right),
    .config_config_addr(Tile_X00_Y0B_config_out_config_addr),
    .config_config_data(Tile_X00_Y0B_config_out_config_data),
    .config_out_config_addr(Tile_X00_Y0C_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y0C_config_out_config_data),
    .config_out_read(Tile_X00_Y0C_config_out_read),
    .config_out_write(Tile_X00_Y0C_config_out_write),
    .config_read(Tile_X00_Y0B_config_out_read),
    .config_write(Tile_X00_Y0B_config_out_write),
    .hi(Tile_X00_Y0C_hi_unq1),
    .lo(Tile_X00_Y0C_lo_unq1),
    .read_config_data(Tile_X00_Y0C_read_config_data),
    .read_config_data_in(Tile_X00_Y0B_read_config_data),
    .reset(Tile_X00_Y0B_reset_out),
    .reset_out(Tile_X00_Y0C_reset_out),
    .stall(Tile_X00_Y0B_stall_out),
    .stall_out(Tile_X00_Y0C_stall_out),
    .tile_id(Tile_X00_Y0C_tile_id_in)
);
mantle_wire__typeBit9 Tile_X00_Y0C_hi (
    .in(Tile_X00_Y0C_hi_unq1),
    .out(Tile_X00_Y0C_hi_out)
);
mantle_wire__typeBit8 Tile_X00_Y0C_lo (
    .in(Tile_X00_Y0C_lo_unq1),
    .out(Tile_X00_Y0C_lo_out)
);
wire [15:0] Tile_X00_Y0C_tile_id_out;
assign Tile_X00_Y0C_tile_id_out = {Tile_X00_Y0C_lo_out[7],Tile_X00_Y0C_lo_out[7:6],Tile_X00_Y0C_lo_out[6:5],Tile_X00_Y0C_lo_out[5:4],Tile_X00_Y0C_lo_out[4:3],Tile_X00_Y0C_lo_out[3:2],Tile_X00_Y0C_lo_out[2],Tile_X00_Y0C_hi_out[2:1],Tile_X00_Y0C_lo_out[0],Tile_X00_Y0C_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X00_Y0C_tile_id (
    .in(Tile_X00_Y0C_tile_id_in),
    .out(Tile_X00_Y0C_tile_id_out)
);
Tile_PE Tile_X00_Y0D (
    .SB_T0_EAST_SB_IN_B1(Tile_X01_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X01_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X00_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X00_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X00_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(const_0_1_out),
    .SB_T0_WEST_SB_IN_B16(const_0_16_out),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X00_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X01_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X01_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X00_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X00_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X00_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(const_0_1_out),
    .SB_T1_WEST_SB_IN_B16(const_0_16_out),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X00_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X01_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X01_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X00_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X00_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X00_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(const_0_1_out),
    .SB_T2_WEST_SB_IN_B16(const_0_16_out),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X00_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X01_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X01_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X00_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X00_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X00_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X00_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X00_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X00_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X00_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(const_0_1_out),
    .SB_T3_WEST_SB_IN_B16(const_0_16_out),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X00_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X01_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X01_Y0D_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X00_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X00_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X00_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X00_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X00_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X00_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X00_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(const_0_1_out),
    .SB_T4_WEST_SB_IN_B16(const_0_16_out),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X00_Y0D_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X00_Y0C_clk_out),
    .clk_out(Tile_X00_Y0D_clk_out),
    .clk_pass_through(Tile_X00_Y0C_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X00_Y0D_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X00_Y0D_clk_pass_through_out_right),
    .config_config_addr(Tile_X00_Y0C_config_out_config_addr),
    .config_config_data(Tile_X00_Y0C_config_out_config_data),
    .config_out_config_addr(Tile_X00_Y0D_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y0D_config_out_config_data),
    .config_out_read(Tile_X00_Y0D_config_out_read),
    .config_out_write(Tile_X00_Y0D_config_out_write),
    .config_read(Tile_X00_Y0C_config_out_read),
    .config_write(Tile_X00_Y0C_config_out_write),
    .hi(Tile_X00_Y0D_hi_unq1),
    .lo(Tile_X00_Y0D_lo_unq1),
    .read_config_data(Tile_X00_Y0D_read_config_data),
    .read_config_data_in(Tile_X00_Y0C_read_config_data),
    .reset(Tile_X00_Y0C_reset_out),
    .reset_out(Tile_X00_Y0D_reset_out),
    .stall(Tile_X00_Y0C_stall_out),
    .stall_out(Tile_X00_Y0D_stall_out),
    .tile_id(Tile_X00_Y0D_tile_id_in)
);
mantle_wire__typeBit9 Tile_X00_Y0D_hi (
    .in(Tile_X00_Y0D_hi_unq1),
    .out(Tile_X00_Y0D_hi_out)
);
mantle_wire__typeBit8 Tile_X00_Y0D_lo (
    .in(Tile_X00_Y0D_lo_unq1),
    .out(Tile_X00_Y0D_lo_out)
);
wire [15:0] Tile_X00_Y0D_tile_id_out;
assign Tile_X00_Y0D_tile_id_out = {Tile_X00_Y0D_lo_out[7],Tile_X00_Y0D_lo_out[7:6],Tile_X00_Y0D_lo_out[6:5],Tile_X00_Y0D_lo_out[5:4],Tile_X00_Y0D_lo_out[4:3],Tile_X00_Y0D_lo_out[3:2],Tile_X00_Y0D_lo_out[2],Tile_X00_Y0D_hi_out[2:1],Tile_X00_Y0D_lo_out[0],Tile_X00_Y0D_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X00_Y0D_tile_id (
    .in(Tile_X00_Y0D_tile_id_in),
    .out(Tile_X00_Y0D_tile_id_out)
);
Tile_PE Tile_X00_Y0E (
    .SB_T0_EAST_SB_IN_B1(Tile_X01_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X01_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X00_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X00_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X00_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(const_0_1_out),
    .SB_T0_WEST_SB_IN_B16(const_0_16_out),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X00_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X01_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X01_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X00_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X00_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X00_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(const_0_1_out),
    .SB_T1_WEST_SB_IN_B16(const_0_16_out),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X00_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X01_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X01_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X00_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X00_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X00_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(const_0_1_out),
    .SB_T2_WEST_SB_IN_B16(const_0_16_out),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X00_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X01_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X01_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X00_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X00_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X00_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X00_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X00_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X00_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X00_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(const_0_1_out),
    .SB_T3_WEST_SB_IN_B16(const_0_16_out),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X00_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X01_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X01_Y0E_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X00_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X00_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X00_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X00_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X00_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X00_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X00_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(const_0_1_out),
    .SB_T4_WEST_SB_IN_B16(const_0_16_out),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X00_Y0E_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X00_Y0D_clk_out),
    .clk_out(Tile_X00_Y0E_clk_out),
    .clk_pass_through(Tile_X00_Y0D_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X00_Y0E_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X00_Y0E_clk_pass_through_out_right),
    .config_config_addr(Tile_X00_Y0D_config_out_config_addr),
    .config_config_data(Tile_X00_Y0D_config_out_config_data),
    .config_out_config_addr(Tile_X00_Y0E_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y0E_config_out_config_data),
    .config_out_read(Tile_X00_Y0E_config_out_read),
    .config_out_write(Tile_X00_Y0E_config_out_write),
    .config_read(Tile_X00_Y0D_config_out_read),
    .config_write(Tile_X00_Y0D_config_out_write),
    .hi(Tile_X00_Y0E_hi_unq1),
    .lo(Tile_X00_Y0E_lo_unq1),
    .read_config_data(Tile_X00_Y0E_read_config_data),
    .read_config_data_in(Tile_X00_Y0D_read_config_data),
    .reset(Tile_X00_Y0D_reset_out),
    .reset_out(Tile_X00_Y0E_reset_out),
    .stall(Tile_X00_Y0D_stall_out),
    .stall_out(Tile_X00_Y0E_stall_out),
    .tile_id(Tile_X00_Y0E_tile_id_in)
);
mantle_wire__typeBit9 Tile_X00_Y0E_hi (
    .in(Tile_X00_Y0E_hi_unq1),
    .out(Tile_X00_Y0E_hi_out)
);
mantle_wire__typeBit8 Tile_X00_Y0E_lo (
    .in(Tile_X00_Y0E_lo_unq1),
    .out(Tile_X00_Y0E_lo_out)
);
wire [15:0] Tile_X00_Y0E_tile_id_out;
assign Tile_X00_Y0E_tile_id_out = {Tile_X00_Y0E_lo_out[7],Tile_X00_Y0E_lo_out[7:6],Tile_X00_Y0E_lo_out[6:5],Tile_X00_Y0E_lo_out[5:4],Tile_X00_Y0E_lo_out[4:3],Tile_X00_Y0E_lo_out[3:2],Tile_X00_Y0E_lo_out[2],Tile_X00_Y0E_hi_out[2:1],Tile_X00_Y0E_hi_out[1],Tile_X00_Y0E_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X00_Y0E_tile_id (
    .in(Tile_X00_Y0E_tile_id_in),
    .out(Tile_X00_Y0E_tile_id_out)
);
Tile_PE Tile_X00_Y0F (
    .SB_T0_EAST_SB_IN_B1(Tile_X01_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X01_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X00_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X00_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X00_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X00_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X00_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(const_0_1_out),
    .SB_T0_WEST_SB_IN_B16(const_0_16_out),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X00_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X01_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X01_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X00_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X00_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X00_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X00_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X00_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(const_0_1_out),
    .SB_T1_WEST_SB_IN_B16(const_0_16_out),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X00_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X01_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X01_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X00_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X00_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X00_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X00_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X00_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(const_0_1_out),
    .SB_T2_WEST_SB_IN_B16(const_0_16_out),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X00_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X01_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X01_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X00_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X00_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X00_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X00_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X00_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X00_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X00_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(const_0_1_out),
    .SB_T3_WEST_SB_IN_B16(const_0_16_out),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X00_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X01_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X01_Y0F_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X00_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X00_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X00_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X00_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X00_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X00_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X00_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(const_0_1_out),
    .SB_T4_WEST_SB_IN_B16(const_0_16_out),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X00_Y0F_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X00_Y0E_clk_out),
    .clk_out(Tile_X00_Y0F_clk_out),
    .clk_pass_through(Tile_X00_Y0E_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X00_Y0F_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X00_Y0F_clk_pass_through_out_right),
    .config_config_addr(Tile_X00_Y0E_config_out_config_addr),
    .config_config_data(Tile_X00_Y0E_config_out_config_data),
    .config_out_config_addr(Tile_X00_Y0F_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y0F_config_out_config_data),
    .config_out_read(Tile_X00_Y0F_config_out_read),
    .config_out_write(Tile_X00_Y0F_config_out_write),
    .config_read(Tile_X00_Y0E_config_out_read),
    .config_write(Tile_X00_Y0E_config_out_write),
    .hi(Tile_X00_Y0F_hi_unq1),
    .lo(Tile_X00_Y0F_lo_unq1),
    .read_config_data(Tile_X00_Y0F_read_config_data),
    .read_config_data_in(Tile_X00_Y0E_read_config_data),
    .reset(Tile_X00_Y0E_reset_out),
    .reset_out(Tile_X00_Y0F_reset_out),
    .stall(Tile_X00_Y0E_stall_out),
    .stall_out(Tile_X00_Y0F_stall_out),
    .tile_id(Tile_X00_Y0F_tile_id_in)
);
mantle_wire__typeBit9 Tile_X00_Y0F_hi (
    .in(Tile_X00_Y0F_hi_unq1),
    .out(Tile_X00_Y0F_hi_out)
);
mantle_wire__typeBit8 Tile_X00_Y0F_lo (
    .in(Tile_X00_Y0F_lo_unq1),
    .out(Tile_X00_Y0F_lo_out)
);
wire [15:0] Tile_X00_Y0F_tile_id_out;
assign Tile_X00_Y0F_tile_id_out = {Tile_X00_Y0F_lo_out[7],Tile_X00_Y0F_lo_out[7:6],Tile_X00_Y0F_lo_out[6:5],Tile_X00_Y0F_lo_out[5:4],Tile_X00_Y0F_lo_out[4:3],Tile_X00_Y0F_lo_out[3:2],Tile_X00_Y0F_lo_out[2],Tile_X00_Y0F_hi_out[2:1],Tile_X00_Y0F_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X00_Y0F_tile_id (
    .in(Tile_X00_Y0F_tile_id_in),
    .out(Tile_X00_Y0F_tile_id_out)
);
Tile_PE Tile_X00_Y10 (
    .SB_T0_EAST_SB_IN_B1(Tile_X01_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X01_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X00_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X00_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X00_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X00_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X00_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X00_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T0_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X00_Y10_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X00_Y10_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(const_0_1_out),
    .SB_T0_WEST_SB_IN_B16(const_0_16_out),
    .SB_T0_WEST_SB_OUT_B1(Tile_X00_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X00_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X01_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X01_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X00_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X00_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X00_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X00_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X00_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X00_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T1_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X00_Y10_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X00_Y10_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(const_0_1_out),
    .SB_T1_WEST_SB_IN_B16(const_0_16_out),
    .SB_T1_WEST_SB_OUT_B1(Tile_X00_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X00_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X01_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X01_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X00_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X00_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X00_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X00_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X00_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X00_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T2_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X00_Y10_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X00_Y10_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(const_0_1_out),
    .SB_T2_WEST_SB_IN_B16(const_0_16_out),
    .SB_T2_WEST_SB_OUT_B1(Tile_X00_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X00_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X01_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X01_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X00_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X00_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X00_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X00_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X00_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X00_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T3_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X00_Y10_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X00_Y10_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(const_0_1_out),
    .SB_T3_WEST_SB_IN_B16(const_0_16_out),
    .SB_T3_WEST_SB_OUT_B1(Tile_X00_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X00_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X01_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X01_Y10_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X00_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X00_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X00_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X00_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X00_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X00_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T4_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X00_Y10_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X00_Y10_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(const_0_1_out),
    .SB_T4_WEST_SB_IN_B16(const_0_16_out),
    .SB_T4_WEST_SB_OUT_B1(Tile_X00_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X00_Y10_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X00_Y0F_clk_out),
    .clk_out(Tile_X00_Y10_clk_out),
    .clk_pass_through(Tile_X00_Y0F_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X00_Y10_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X00_Y10_clk_pass_through_out_right),
    .config_config_addr(Tile_X00_Y0F_config_out_config_addr),
    .config_config_data(Tile_X00_Y0F_config_out_config_data),
    .config_out_config_addr(Tile_X00_Y10_config_out_config_addr),
    .config_out_config_data(Tile_X00_Y10_config_out_config_data),
    .config_out_read(Tile_X00_Y10_config_out_read),
    .config_out_write(Tile_X00_Y10_config_out_write),
    .config_read(Tile_X00_Y0F_config_out_read),
    .config_write(Tile_X00_Y0F_config_out_write),
    .hi(Tile_X00_Y10_hi),
    .lo(Tile_X00_Y10_lo_unq1),
    .read_config_data(Tile_X00_Y10_read_config_data),
    .read_config_data_in(Tile_X00_Y0F_read_config_data),
    .reset(Tile_X00_Y0F_reset_out),
    .reset_out(Tile_X00_Y10_reset_out),
    .stall(Tile_X00_Y0F_stall_out),
    .stall_out(Tile_X00_Y10_stall_out),
    .tile_id(Tile_X00_Y10_tile_id_in)
);
mantle_wire__typeBit8 Tile_X00_Y10_lo (
    .in(Tile_X00_Y10_lo_unq1),
    .out(Tile_X00_Y10_lo_out)
);
wire [15:0] Tile_X00_Y10_tile_id_out;
assign Tile_X00_Y10_tile_id_out = {Tile_X00_Y10_lo_out[7],Tile_X00_Y10_lo_out[7:6],Tile_X00_Y10_lo_out[6:5],Tile_X00_Y10_lo_out[5:4],Tile_X00_Y10_lo_out[4:3],Tile_X00_Y10_lo_out[3:2],Tile_X00_Y10_hi[2],Tile_X00_Y10_lo_out[1],Tile_X00_Y10_lo_out[1:0],Tile_X00_Y10_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X00_Y10_tile_id (
    .in(Tile_X00_Y10_tile_id_in),
    .out(Tile_X00_Y10_tile_id_out)
);
wire [15:0] Tile_X01_Y00_tile_id;
assign Tile_X01_Y00_tile_id = {Tile_X01_Y00_lo[7],Tile_X01_Y00_lo[7:6],Tile_X01_Y00_lo[6:5],Tile_X01_Y00_lo[5:4],Tile_X01_Y00_hi[4],Tile_X01_Y00_lo[3],Tile_X01_Y00_lo[3:2],Tile_X01_Y00_lo[2:1],Tile_X01_Y00_lo[1:0],Tile_X01_Y00_lo[0]};
Tile_io_core Tile_X01_Y00 (
    .tile_id(Tile_X01_Y00_tile_id),
    .glb2io_1(glb2io_1_X01_Y00),
    .f2io_1(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B1),
    .io2glb_1(Tile_X01_Y00_io2glb_1),
    .io2f_1(Tile_X01_Y00_io2f_1),
    .glb2io_16(glb2io_16_X01_Y00),
    .f2io_16(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B16),
    .io2glb_16(Tile_X01_Y00_io2glb_16),
    .io2f_16(Tile_X01_Y00_io2f_16),
    .hi(Tile_X01_Y00_hi),
    .lo(Tile_X01_Y00_lo)
);
Tile_PE Tile_X01_Y01 (
    .SB_T0_EAST_SB_IN_B1(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X01_Y00_io2f_1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X01_Y00_io2f_16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y01_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X00_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X01_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X01_Y00_io2f_1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X01_Y00_io2f_16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y01_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X00_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X01_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X01_Y00_io2f_1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X01_Y00_io2f_16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y01_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X00_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X01_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X02_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X02_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X01_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X01_Y00_io2f_1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X01_Y00_io2f_16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y01_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X01_Y01_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X00_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X00_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X01_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X02_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X02_Y01_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X01_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X01_Y00_io2f_1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X01_Y00_io2f_16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y01_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X01_Y01_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X00_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X00_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X01_Y01_SB_T4_WEST_SB_OUT_B16),
    .clk(clk),
    .clk_out(Tile_X01_Y01_clk_out),
    .clk_pass_through(clk),
    .clk_pass_through_out_bot(Tile_X01_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X01_Y01_clk_pass_through_out_right),
    .config_config_addr(config_1_config_addr),
    .config_config_data(config_1_config_data),
    .config_out_config_addr(Tile_X01_Y01_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y01_config_out_config_data),
    .config_out_read(Tile_X01_Y01_config_out_read),
    .config_out_write(Tile_X01_Y01_config_out_write),
    .config_read(config_1_read),
    .config_write(config_1_write),
    .hi(Tile_X01_Y01_hi),
    .lo(Tile_X01_Y01_lo_unq1),
    .read_config_data(Tile_X01_Y01_read_config_data),
    .read_config_data_in(const_0_32_out),
    .reset(reset),
    .reset_out(Tile_X01_Y01_reset_out),
    .stall(stall[1]),
    .stall_out(Tile_X01_Y01_stall_out),
    .tile_id(Tile_X01_Y01_tile_id_in)
);
mantle_wire__typeBit8 Tile_X01_Y01_lo (
    .in(Tile_X01_Y01_lo_unq1),
    .out(Tile_X01_Y01_lo_out)
);
wire [15:0] Tile_X01_Y01_tile_id_out;
assign Tile_X01_Y01_tile_id_out = {Tile_X01_Y01_lo_out[7],Tile_X01_Y01_lo_out[7:6],Tile_X01_Y01_lo_out[6:5],Tile_X01_Y01_lo_out[5:4],Tile_X01_Y01_hi[4],Tile_X01_Y01_lo_out[3],Tile_X01_Y01_lo_out[3:2],Tile_X01_Y01_lo_out[2:1],Tile_X01_Y01_lo_out[1:0],Tile_X01_Y01_hi[0]};
mantle_wire__typeBitIn16 Tile_X01_Y01_tile_id (
    .in(Tile_X01_Y01_tile_id_in),
    .out(Tile_X01_Y01_tile_id_out)
);
Tile_PE Tile_X01_Y02 (
    .SB_T0_EAST_SB_IN_B1(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X01_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X00_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X01_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X01_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X00_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X01_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X01_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X00_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X01_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X02_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X02_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X01_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X01_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X01_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X00_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X00_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X01_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X02_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X02_Y02_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X01_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X01_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X01_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X00_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X00_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X01_Y02_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X01_Y01_clk_out),
    .clk_out(Tile_X01_Y02_clk_out),
    .clk_pass_through(Tile_X01_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X01_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X01_Y02_clk_pass_through_out_right),
    .config_config_addr(Tile_X01_Y01_config_out_config_addr),
    .config_config_data(Tile_X01_Y01_config_out_config_data),
    .config_out_config_addr(Tile_X01_Y02_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y02_config_out_config_data),
    .config_out_read(Tile_X01_Y02_config_out_read),
    .config_out_write(Tile_X01_Y02_config_out_write),
    .config_read(Tile_X01_Y01_config_out_read),
    .config_write(Tile_X01_Y01_config_out_write),
    .hi(Tile_X01_Y02_hi),
    .lo(Tile_X01_Y02_lo_unq1),
    .read_config_data(Tile_X01_Y02_read_config_data),
    .read_config_data_in(Tile_X01_Y01_read_config_data),
    .reset(Tile_X01_Y01_reset_out),
    .reset_out(Tile_X01_Y02_reset_out),
    .stall(Tile_X01_Y01_stall_out),
    .stall_out(Tile_X01_Y02_stall_out),
    .tile_id(Tile_X01_Y02_tile_id_in)
);
mantle_wire__typeBit8 Tile_X01_Y02_lo (
    .in(Tile_X01_Y02_lo_unq1),
    .out(Tile_X01_Y02_lo_out)
);
wire [15:0] Tile_X01_Y02_tile_id_out;
assign Tile_X01_Y02_tile_id_out = {Tile_X01_Y02_lo_out[7],Tile_X01_Y02_lo_out[7:6],Tile_X01_Y02_lo_out[6:5],Tile_X01_Y02_lo_out[5:4],Tile_X01_Y02_hi[4],Tile_X01_Y02_lo_out[3],Tile_X01_Y02_lo_out[3:2],Tile_X01_Y02_lo_out[2:1],Tile_X01_Y02_lo_out[1],Tile_X01_Y02_hi[1],Tile_X01_Y02_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X01_Y02_tile_id (
    .in(Tile_X01_Y02_tile_id_in),
    .out(Tile_X01_Y02_tile_id_out)
);
Tile_PE Tile_X01_Y03 (
    .SB_T0_EAST_SB_IN_B1(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X01_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X00_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X01_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X01_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X00_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X01_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X01_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X00_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X01_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X02_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X02_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X01_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X01_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X01_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X00_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X00_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X01_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X02_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X02_Y03_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X01_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X01_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X01_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X00_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X00_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X01_Y03_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X01_Y02_clk_out),
    .clk_out(Tile_X01_Y03_clk_out),
    .clk_pass_through(Tile_X01_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X01_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X01_Y03_clk_pass_through_out_right),
    .config_config_addr(Tile_X01_Y02_config_out_config_addr),
    .config_config_data(Tile_X01_Y02_config_out_config_data),
    .config_out_config_addr(Tile_X01_Y03_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y03_config_out_config_data),
    .config_out_read(Tile_X01_Y03_config_out_read),
    .config_out_write(Tile_X01_Y03_config_out_write),
    .config_read(Tile_X01_Y02_config_out_read),
    .config_write(Tile_X01_Y02_config_out_write),
    .hi(Tile_X01_Y03_hi_unq1),
    .lo(Tile_X01_Y03_lo_unq1),
    .read_config_data(Tile_X01_Y03_read_config_data),
    .read_config_data_in(Tile_X01_Y02_read_config_data),
    .reset(Tile_X01_Y02_reset_out),
    .reset_out(Tile_X01_Y03_reset_out),
    .stall(Tile_X01_Y02_stall_out),
    .stall_out(Tile_X01_Y03_stall_out),
    .tile_id(Tile_X01_Y03_tile_id_in)
);
mantle_wire__typeBit9 Tile_X01_Y03_hi (
    .in(Tile_X01_Y03_hi_unq1),
    .out(Tile_X01_Y03_hi_out)
);
mantle_wire__typeBit8 Tile_X01_Y03_lo (
    .in(Tile_X01_Y03_lo_unq1),
    .out(Tile_X01_Y03_lo_out)
);
wire [15:0] Tile_X01_Y03_tile_id_out;
assign Tile_X01_Y03_tile_id_out = {Tile_X01_Y03_lo_out[7],Tile_X01_Y03_lo_out[7:6],Tile_X01_Y03_lo_out[6:5],Tile_X01_Y03_lo_out[5:4],Tile_X01_Y03_hi_out[4],Tile_X01_Y03_lo_out[3],Tile_X01_Y03_lo_out[3:2],Tile_X01_Y03_lo_out[2:1],Tile_X01_Y03_lo_out[1],Tile_X01_Y03_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X01_Y03_tile_id (
    .in(Tile_X01_Y03_tile_id_in),
    .out(Tile_X01_Y03_tile_id_out)
);
Tile_PE Tile_X01_Y04 (
    .SB_T0_EAST_SB_IN_B1(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X01_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X00_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X01_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X01_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X00_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X01_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X01_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X00_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X01_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X02_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X02_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X01_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X01_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X01_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X01_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X01_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X00_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X00_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X01_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X02_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X02_Y04_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X01_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X01_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X01_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X01_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X01_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X00_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X00_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X01_Y04_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X01_Y03_clk_out),
    .clk_out(Tile_X01_Y04_clk_out),
    .clk_pass_through(Tile_X01_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X01_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X01_Y04_clk_pass_through_out_right),
    .config_config_addr(Tile_X01_Y03_config_out_config_addr),
    .config_config_data(Tile_X01_Y03_config_out_config_data),
    .config_out_config_addr(Tile_X01_Y04_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y04_config_out_config_data),
    .config_out_read(Tile_X01_Y04_config_out_read),
    .config_out_write(Tile_X01_Y04_config_out_write),
    .config_read(Tile_X01_Y03_config_out_read),
    .config_write(Tile_X01_Y03_config_out_write),
    .hi(Tile_X01_Y04_hi),
    .lo(Tile_X01_Y04_lo_unq1),
    .read_config_data(Tile_X01_Y04_read_config_data),
    .read_config_data_in(Tile_X01_Y03_read_config_data),
    .reset(Tile_X01_Y03_reset_out),
    .reset_out(Tile_X01_Y04_reset_out),
    .stall(Tile_X01_Y03_stall_out),
    .stall_out(Tile_X01_Y04_stall_out),
    .tile_id(Tile_X01_Y04_tile_id_in)
);
mantle_wire__typeBit8 Tile_X01_Y04_lo (
    .in(Tile_X01_Y04_lo_unq1),
    .out(Tile_X01_Y04_lo_out)
);
wire [15:0] Tile_X01_Y04_tile_id_out;
assign Tile_X01_Y04_tile_id_out = {Tile_X01_Y04_lo_out[7],Tile_X01_Y04_lo_out[7:6],Tile_X01_Y04_lo_out[6:5],Tile_X01_Y04_lo_out[5:4],Tile_X01_Y04_hi[4],Tile_X01_Y04_lo_out[3],Tile_X01_Y04_lo_out[3:2],Tile_X01_Y04_lo_out[2:1],Tile_X01_Y04_hi[1],Tile_X01_Y04_lo_out[0],Tile_X01_Y04_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X01_Y04_tile_id (
    .in(Tile_X01_Y04_tile_id_in),
    .out(Tile_X01_Y04_tile_id_out)
);
Tile_PE Tile_X01_Y05 (
    .SB_T0_EAST_SB_IN_B1(Tile_X02_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X02_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X01_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X01_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X00_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X00_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X01_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X02_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X02_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X01_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X01_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X00_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X00_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X01_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X02_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X02_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X01_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X01_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X00_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X00_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X01_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X02_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X02_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X01_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X01_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X01_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X01_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X01_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X01_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X00_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X00_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X01_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X02_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X02_Y05_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X01_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X01_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X01_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X01_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X01_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X01_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X00_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X00_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X01_Y05_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X01_Y04_clk_out),
    .clk_out(Tile_X01_Y05_clk_out),
    .clk_pass_through(Tile_X01_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X01_Y05_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X01_Y05_clk_pass_through_out_right),
    .config_config_addr(Tile_X01_Y04_config_out_config_addr),
    .config_config_data(Tile_X01_Y04_config_out_config_data),
    .config_out_config_addr(Tile_X01_Y05_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y05_config_out_config_data),
    .config_out_read(Tile_X01_Y05_config_out_read),
    .config_out_write(Tile_X01_Y05_config_out_write),
    .config_read(Tile_X01_Y04_config_out_read),
    .config_write(Tile_X01_Y04_config_out_write),
    .hi(Tile_X01_Y05_hi),
    .lo(Tile_X01_Y05_lo_unq1),
    .read_config_data(Tile_X01_Y05_read_config_data),
    .read_config_data_in(Tile_X01_Y04_read_config_data),
    .reset(Tile_X01_Y04_reset_out),
    .reset_out(Tile_X01_Y05_reset_out),
    .stall(Tile_X01_Y04_stall_out),
    .stall_out(Tile_X01_Y05_stall_out),
    .tile_id(Tile_X01_Y05_tile_id_in)
);
mantle_wire__typeBit8 Tile_X01_Y05_lo (
    .in(Tile_X01_Y05_lo_unq1),
    .out(Tile_X01_Y05_lo_out)
);
wire [15:0] Tile_X01_Y05_tile_id_out;
assign Tile_X01_Y05_tile_id_out = {Tile_X01_Y05_lo_out[7],Tile_X01_Y05_lo_out[7:6],Tile_X01_Y05_lo_out[6:5],Tile_X01_Y05_lo_out[5:4],Tile_X01_Y05_hi[4],Tile_X01_Y05_lo_out[3],Tile_X01_Y05_lo_out[3:2],Tile_X01_Y05_lo_out[2:1],Tile_X01_Y05_hi[1],Tile_X01_Y05_lo_out[0],Tile_X01_Y05_hi[0]};
mantle_wire__typeBitIn16 Tile_X01_Y05_tile_id (
    .in(Tile_X01_Y05_tile_id_in),
    .out(Tile_X01_Y05_tile_id_out)
);
Tile_PE Tile_X01_Y06 (
    .SB_T0_EAST_SB_IN_B1(Tile_X02_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X02_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X01_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X01_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X01_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X00_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X00_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X01_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X02_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X02_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X01_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X01_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X01_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X00_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X00_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X01_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X02_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X02_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X01_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X01_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X01_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X00_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X00_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X01_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X02_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X02_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X01_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X01_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X01_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X01_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X01_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X01_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X01_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X00_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X00_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X01_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X02_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X02_Y06_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X01_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X01_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X01_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X01_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X01_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X01_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X01_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X00_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X00_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X01_Y06_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X01_Y05_clk_out),
    .clk_out(Tile_X01_Y06_clk_out),
    .clk_pass_through(Tile_X01_Y05_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X01_Y06_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X01_Y06_clk_pass_through_out_right),
    .config_config_addr(Tile_X01_Y05_config_out_config_addr),
    .config_config_data(Tile_X01_Y05_config_out_config_data),
    .config_out_config_addr(Tile_X01_Y06_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y06_config_out_config_data),
    .config_out_read(Tile_X01_Y06_config_out_read),
    .config_out_write(Tile_X01_Y06_config_out_write),
    .config_read(Tile_X01_Y05_config_out_read),
    .config_write(Tile_X01_Y05_config_out_write),
    .hi(Tile_X01_Y06_hi),
    .lo(Tile_X01_Y06_lo_unq1),
    .read_config_data(Tile_X01_Y06_read_config_data),
    .read_config_data_in(Tile_X01_Y05_read_config_data),
    .reset(Tile_X01_Y05_reset_out),
    .reset_out(Tile_X01_Y06_reset_out),
    .stall(Tile_X01_Y05_stall_out),
    .stall_out(Tile_X01_Y06_stall_out),
    .tile_id(Tile_X01_Y06_tile_id_in)
);
mantle_wire__typeBit8 Tile_X01_Y06_lo (
    .in(Tile_X01_Y06_lo_unq1),
    .out(Tile_X01_Y06_lo_out)
);
wire [15:0] Tile_X01_Y06_tile_id_out;
assign Tile_X01_Y06_tile_id_out = {Tile_X01_Y06_lo_out[7],Tile_X01_Y06_lo_out[7:6],Tile_X01_Y06_lo_out[6:5],Tile_X01_Y06_lo_out[5:4],Tile_X01_Y06_hi[4],Tile_X01_Y06_lo_out[3],Tile_X01_Y06_lo_out[3:2],Tile_X01_Y06_lo_out[2:1],Tile_X01_Y06_hi[1],Tile_X01_Y06_hi[1],Tile_X01_Y06_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X01_Y06_tile_id (
    .in(Tile_X01_Y06_tile_id_in),
    .out(Tile_X01_Y06_tile_id_out)
);
Tile_PE Tile_X01_Y07 (
    .SB_T0_EAST_SB_IN_B1(Tile_X02_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X02_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X01_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X01_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X01_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X00_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X00_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X01_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X02_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X02_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X01_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X01_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X01_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X00_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X00_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X01_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X02_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X02_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X01_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X01_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X01_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X00_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X00_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X01_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X02_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X02_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X01_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X01_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X01_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X01_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X01_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X01_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X01_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X00_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X00_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X01_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X02_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X02_Y07_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X01_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X01_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X01_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X01_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X01_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X01_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X01_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X00_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X00_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X01_Y07_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X01_Y06_clk_out),
    .clk_out(Tile_X01_Y07_clk_out),
    .clk_pass_through(Tile_X01_Y06_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X01_Y07_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X01_Y07_clk_pass_through_out_right),
    .config_config_addr(Tile_X01_Y06_config_out_config_addr),
    .config_config_data(Tile_X01_Y06_config_out_config_data),
    .config_out_config_addr(Tile_X01_Y07_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y07_config_out_config_data),
    .config_out_read(Tile_X01_Y07_config_out_read),
    .config_out_write(Tile_X01_Y07_config_out_write),
    .config_read(Tile_X01_Y06_config_out_read),
    .config_write(Tile_X01_Y06_config_out_write),
    .hi(Tile_X01_Y07_hi_unq1),
    .lo(Tile_X01_Y07_lo_unq1),
    .read_config_data(Tile_X01_Y07_read_config_data),
    .read_config_data_in(Tile_X01_Y06_read_config_data),
    .reset(Tile_X01_Y06_reset_out),
    .reset_out(Tile_X01_Y07_reset_out),
    .stall(Tile_X01_Y06_stall_out),
    .stall_out(Tile_X01_Y07_stall_out),
    .tile_id(Tile_X01_Y07_tile_id_in)
);
mantle_wire__typeBit9 Tile_X01_Y07_hi (
    .in(Tile_X01_Y07_hi_unq1),
    .out(Tile_X01_Y07_hi_out)
);
mantle_wire__typeBit8 Tile_X01_Y07_lo (
    .in(Tile_X01_Y07_lo_unq1),
    .out(Tile_X01_Y07_lo_out)
);
wire [15:0] Tile_X01_Y07_tile_id_out;
assign Tile_X01_Y07_tile_id_out = {Tile_X01_Y07_lo_out[7],Tile_X01_Y07_lo_out[7:6],Tile_X01_Y07_lo_out[6:5],Tile_X01_Y07_lo_out[5:4],Tile_X01_Y07_hi_out[4],Tile_X01_Y07_lo_out[3],Tile_X01_Y07_lo_out[3:2],Tile_X01_Y07_lo_out[2:1],Tile_X01_Y07_hi_out[1],Tile_X01_Y07_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X01_Y07_tile_id (
    .in(Tile_X01_Y07_tile_id_in),
    .out(Tile_X01_Y07_tile_id_out)
);
Tile_PE Tile_X01_Y08 (
    .SB_T0_EAST_SB_IN_B1(Tile_X02_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X02_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X01_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X01_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X01_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X00_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X00_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X01_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X02_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X02_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X01_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X01_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X01_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X00_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X00_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X01_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X02_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X02_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X01_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X01_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X01_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X00_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X00_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X01_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X02_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X02_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X01_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X01_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X01_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X01_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X01_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X01_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X01_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X00_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X00_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X01_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X02_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X02_Y08_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X01_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X01_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X01_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X01_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X01_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X01_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X01_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X00_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X00_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X01_Y08_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X01_Y07_clk_out),
    .clk_out(Tile_X01_Y08_clk_out),
    .clk_pass_through(Tile_X01_Y07_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X01_Y08_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X01_Y08_clk_pass_through_out_right),
    .config_config_addr(Tile_X01_Y07_config_out_config_addr),
    .config_config_data(Tile_X01_Y07_config_out_config_data),
    .config_out_config_addr(Tile_X01_Y08_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y08_config_out_config_data),
    .config_out_read(Tile_X01_Y08_config_out_read),
    .config_out_write(Tile_X01_Y08_config_out_write),
    .config_read(Tile_X01_Y07_config_out_read),
    .config_write(Tile_X01_Y07_config_out_write),
    .hi(Tile_X01_Y08_hi),
    .lo(Tile_X01_Y08_lo_unq1),
    .read_config_data(Tile_X01_Y08_read_config_data),
    .read_config_data_in(Tile_X01_Y07_read_config_data),
    .reset(Tile_X01_Y07_reset_out),
    .reset_out(Tile_X01_Y08_reset_out),
    .stall(Tile_X01_Y07_stall_out),
    .stall_out(Tile_X01_Y08_stall_out),
    .tile_id(Tile_X01_Y08_tile_id_in)
);
mantle_wire__typeBit8 Tile_X01_Y08_lo (
    .in(Tile_X01_Y08_lo_unq1),
    .out(Tile_X01_Y08_lo_out)
);
wire [15:0] Tile_X01_Y08_tile_id_out;
assign Tile_X01_Y08_tile_id_out = {Tile_X01_Y08_lo_out[7],Tile_X01_Y08_lo_out[7:6],Tile_X01_Y08_lo_out[6:5],Tile_X01_Y08_lo_out[5:4],Tile_X01_Y08_hi[4],Tile_X01_Y08_lo_out[3],Tile_X01_Y08_lo_out[3:2],Tile_X01_Y08_lo_out[2],Tile_X01_Y08_hi[2],Tile_X01_Y08_lo_out[1:0],Tile_X01_Y08_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X01_Y08_tile_id (
    .in(Tile_X01_Y08_tile_id_in),
    .out(Tile_X01_Y08_tile_id_out)
);
Tile_PE Tile_X01_Y09 (
    .SB_T0_EAST_SB_IN_B1(Tile_X02_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X02_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X01_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X01_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X01_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X00_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X00_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X01_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X02_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X02_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X01_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X01_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X01_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X00_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X00_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X01_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X02_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X02_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X01_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X01_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X01_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X00_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X00_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X01_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X02_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X02_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X01_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X01_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X01_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X01_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X01_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X01_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X01_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X00_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X00_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X01_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X02_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X02_Y09_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X01_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X01_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X01_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X01_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X01_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X01_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X01_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X00_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X00_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X01_Y09_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X01_Y08_clk_out),
    .clk_out(Tile_X01_Y09_clk_out),
    .clk_pass_through(Tile_X01_Y08_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X01_Y09_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X01_Y09_clk_pass_through_out_right),
    .config_config_addr(ConfigPipeStage_inst1_config_out_config_addr),
    .config_config_data(ConfigPipeStage_inst1_config_out_config_data),
    .config_out_config_addr(Tile_X01_Y09_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y09_config_out_config_data),
    .config_out_read(Tile_X01_Y09_config_out_read),
    .config_out_write(Tile_X01_Y09_config_out_write),
    .config_read(ConfigPipeStage_inst1_config_out_read),
    .config_write(ConfigPipeStage_inst1_config_out_write),
    .hi(Tile_X01_Y09_hi),
    .lo(Tile_X01_Y09_lo_unq1),
    .read_config_data(Tile_X01_Y09_read_config_data),
    .read_config_data_in(Tile_X01_Y08_read_config_data),
    .reset(Tile_X01_Y08_reset_out),
    .reset_out(Tile_X01_Y09_reset_out),
    .stall(Tile_X01_Y08_stall_out),
    .stall_out(Tile_X01_Y09_stall_out),
    .tile_id(Tile_X01_Y09_tile_id_in)
);
mantle_wire__typeBit8 Tile_X01_Y09_lo (
    .in(Tile_X01_Y09_lo_unq1),
    .out(Tile_X01_Y09_lo_out)
);
wire [15:0] Tile_X01_Y09_tile_id_out;
assign Tile_X01_Y09_tile_id_out = {Tile_X01_Y09_lo_out[7],Tile_X01_Y09_lo_out[7:6],Tile_X01_Y09_lo_out[6:5],Tile_X01_Y09_lo_out[5:4],Tile_X01_Y09_hi[4],Tile_X01_Y09_lo_out[3],Tile_X01_Y09_lo_out[3:2],Tile_X01_Y09_lo_out[2],Tile_X01_Y09_hi[2],Tile_X01_Y09_lo_out[1:0],Tile_X01_Y09_hi[0]};
mantle_wire__typeBitIn16 Tile_X01_Y09_tile_id (
    .in(Tile_X01_Y09_tile_id_in),
    .out(Tile_X01_Y09_tile_id_out)
);
Tile_PE Tile_X01_Y0A (
    .SB_T0_EAST_SB_IN_B1(Tile_X02_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X02_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X01_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X01_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X01_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X00_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X00_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X01_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X02_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X02_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X01_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X01_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X01_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X00_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X00_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X01_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X02_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X02_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X01_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X01_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X01_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X00_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X00_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X01_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X02_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X02_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X01_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X01_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X01_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X01_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X01_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X01_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X01_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X00_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X00_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X01_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X02_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X02_Y0A_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X01_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X01_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X01_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X01_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X01_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X01_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X01_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X00_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X00_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X01_Y0A_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X01_Y09_clk_out),
    .clk_out(Tile_X01_Y0A_clk_out),
    .clk_pass_through(Tile_X01_Y09_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X01_Y0A_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X01_Y0A_clk_pass_through_out_right),
    .config_config_addr(Tile_X01_Y09_config_out_config_addr),
    .config_config_data(Tile_X01_Y09_config_out_config_data),
    .config_out_config_addr(Tile_X01_Y0A_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y0A_config_out_config_data),
    .config_out_read(Tile_X01_Y0A_config_out_read),
    .config_out_write(Tile_X01_Y0A_config_out_write),
    .config_read(Tile_X01_Y09_config_out_read),
    .config_write(Tile_X01_Y09_config_out_write),
    .hi(Tile_X01_Y0A_hi),
    .lo(Tile_X01_Y0A_lo_unq1),
    .read_config_data(Tile_X01_Y0A_read_config_data),
    .read_config_data_in(Tile_X01_Y09_read_config_data),
    .reset(Tile_X01_Y09_reset_out),
    .reset_out(Tile_X01_Y0A_reset_out),
    .stall(Tile_X01_Y09_stall_out),
    .stall_out(Tile_X01_Y0A_stall_out),
    .tile_id(Tile_X01_Y0A_tile_id_in)
);
mantle_wire__typeBit8 Tile_X01_Y0A_lo (
    .in(Tile_X01_Y0A_lo_unq1),
    .out(Tile_X01_Y0A_lo_out)
);
wire [15:0] Tile_X01_Y0A_tile_id_out;
assign Tile_X01_Y0A_tile_id_out = {Tile_X01_Y0A_lo_out[7],Tile_X01_Y0A_lo_out[7:6],Tile_X01_Y0A_lo_out[6:5],Tile_X01_Y0A_lo_out[5:4],Tile_X01_Y0A_hi[4],Tile_X01_Y0A_lo_out[3],Tile_X01_Y0A_lo_out[3:2],Tile_X01_Y0A_lo_out[2],Tile_X01_Y0A_hi[2],Tile_X01_Y0A_lo_out[1],Tile_X01_Y0A_hi[1],Tile_X01_Y0A_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X01_Y0A_tile_id (
    .in(Tile_X01_Y0A_tile_id_in),
    .out(Tile_X01_Y0A_tile_id_out)
);
Tile_PE Tile_X01_Y0B (
    .SB_T0_EAST_SB_IN_B1(Tile_X02_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X02_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X01_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X01_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X01_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X00_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X00_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X01_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X02_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X02_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X01_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X01_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X01_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X00_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X00_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X01_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X02_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X02_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X01_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X01_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X01_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X00_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X00_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X01_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X02_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X02_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X01_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X01_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X01_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X01_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X01_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X01_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X01_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X00_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X00_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X01_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X02_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X02_Y0B_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X01_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X01_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X01_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X01_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X01_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X01_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X01_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X00_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X00_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X01_Y0B_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X01_Y0A_clk_out),
    .clk_out(Tile_X01_Y0B_clk_out),
    .clk_pass_through(Tile_X01_Y0A_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X01_Y0B_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X01_Y0B_clk_pass_through_out_right),
    .config_config_addr(Tile_X01_Y0A_config_out_config_addr),
    .config_config_data(Tile_X01_Y0A_config_out_config_data),
    .config_out_config_addr(Tile_X01_Y0B_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y0B_config_out_config_data),
    .config_out_read(Tile_X01_Y0B_config_out_read),
    .config_out_write(Tile_X01_Y0B_config_out_write),
    .config_read(Tile_X01_Y0A_config_out_read),
    .config_write(Tile_X01_Y0A_config_out_write),
    .hi(Tile_X01_Y0B_hi_unq1),
    .lo(Tile_X01_Y0B_lo_unq1),
    .read_config_data(Tile_X01_Y0B_read_config_data),
    .read_config_data_in(Tile_X01_Y0A_read_config_data),
    .reset(Tile_X01_Y0A_reset_out),
    .reset_out(Tile_X01_Y0B_reset_out),
    .stall(Tile_X01_Y0A_stall_out),
    .stall_out(Tile_X01_Y0B_stall_out),
    .tile_id(Tile_X01_Y0B_tile_id_in)
);
mantle_wire__typeBit9 Tile_X01_Y0B_hi (
    .in(Tile_X01_Y0B_hi_unq1),
    .out(Tile_X01_Y0B_hi_out)
);
mantle_wire__typeBit8 Tile_X01_Y0B_lo (
    .in(Tile_X01_Y0B_lo_unq1),
    .out(Tile_X01_Y0B_lo_out)
);
wire [15:0] Tile_X01_Y0B_tile_id_out;
assign Tile_X01_Y0B_tile_id_out = {Tile_X01_Y0B_lo_out[7],Tile_X01_Y0B_lo_out[7:6],Tile_X01_Y0B_lo_out[6:5],Tile_X01_Y0B_lo_out[5:4],Tile_X01_Y0B_hi_out[4],Tile_X01_Y0B_lo_out[3],Tile_X01_Y0B_lo_out[3:2],Tile_X01_Y0B_lo_out[2],Tile_X01_Y0B_hi_out[2],Tile_X01_Y0B_lo_out[1],Tile_X01_Y0B_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X01_Y0B_tile_id (
    .in(Tile_X01_Y0B_tile_id_in),
    .out(Tile_X01_Y0B_tile_id_out)
);
Tile_PE Tile_X01_Y0C (
    .SB_T0_EAST_SB_IN_B1(Tile_X02_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X02_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X01_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X01_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X01_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X00_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X00_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X01_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X02_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X02_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X01_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X01_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X01_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X00_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X00_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X01_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X02_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X02_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X01_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X01_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X01_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X00_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X00_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X01_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X02_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X02_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X01_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X01_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X01_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X01_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X01_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X01_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X01_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X00_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X00_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X01_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X02_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X02_Y0C_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X01_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X01_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X01_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X01_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X01_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X01_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X01_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X00_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X00_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X01_Y0C_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X01_Y0B_clk_out),
    .clk_out(Tile_X01_Y0C_clk_out),
    .clk_pass_through(Tile_X01_Y0B_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X01_Y0C_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X01_Y0C_clk_pass_through_out_right),
    .config_config_addr(Tile_X01_Y0B_config_out_config_addr),
    .config_config_data(Tile_X01_Y0B_config_out_config_data),
    .config_out_config_addr(Tile_X01_Y0C_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y0C_config_out_config_data),
    .config_out_read(Tile_X01_Y0C_config_out_read),
    .config_out_write(Tile_X01_Y0C_config_out_write),
    .config_read(Tile_X01_Y0B_config_out_read),
    .config_write(Tile_X01_Y0B_config_out_write),
    .hi(Tile_X01_Y0C_hi_unq1),
    .lo(Tile_X01_Y0C_lo_unq1),
    .read_config_data(Tile_X01_Y0C_read_config_data),
    .read_config_data_in(Tile_X01_Y0B_read_config_data),
    .reset(Tile_X01_Y0B_reset_out),
    .reset_out(Tile_X01_Y0C_reset_out),
    .stall(Tile_X01_Y0B_stall_out),
    .stall_out(Tile_X01_Y0C_stall_out),
    .tile_id(Tile_X01_Y0C_tile_id_in)
);
mantle_wire__typeBit9 Tile_X01_Y0C_hi (
    .in(Tile_X01_Y0C_hi_unq1),
    .out(Tile_X01_Y0C_hi_out)
);
mantle_wire__typeBit8 Tile_X01_Y0C_lo (
    .in(Tile_X01_Y0C_lo_unq1),
    .out(Tile_X01_Y0C_lo_out)
);
wire [15:0] Tile_X01_Y0C_tile_id_out;
assign Tile_X01_Y0C_tile_id_out = {Tile_X01_Y0C_lo_out[7],Tile_X01_Y0C_lo_out[7:6],Tile_X01_Y0C_lo_out[6:5],Tile_X01_Y0C_lo_out[5:4],Tile_X01_Y0C_hi_out[4],Tile_X01_Y0C_lo_out[3],Tile_X01_Y0C_lo_out[3:2],Tile_X01_Y0C_lo_out[2],Tile_X01_Y0C_hi_out[2:1],Tile_X01_Y0C_lo_out[0],Tile_X01_Y0C_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X01_Y0C_tile_id (
    .in(Tile_X01_Y0C_tile_id_in),
    .out(Tile_X01_Y0C_tile_id_out)
);
Tile_PE Tile_X01_Y0D (
    .SB_T0_EAST_SB_IN_B1(Tile_X02_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X02_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X01_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X01_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X01_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X00_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X00_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X01_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X02_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X02_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X01_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X01_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X01_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X00_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X00_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X01_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X02_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X02_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X01_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X01_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X01_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X00_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X00_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X01_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X02_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X02_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X01_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X01_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X01_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X01_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X01_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X01_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X01_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X00_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X00_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X01_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X02_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X02_Y0D_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X01_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X01_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X01_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X01_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X01_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X01_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X01_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X00_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X00_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X01_Y0D_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X01_Y0C_clk_out),
    .clk_out(Tile_X01_Y0D_clk_out),
    .clk_pass_through(Tile_X01_Y0C_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X01_Y0D_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X01_Y0D_clk_pass_through_out_right),
    .config_config_addr(Tile_X01_Y0C_config_out_config_addr),
    .config_config_data(Tile_X01_Y0C_config_out_config_data),
    .config_out_config_addr(Tile_X01_Y0D_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y0D_config_out_config_data),
    .config_out_read(Tile_X01_Y0D_config_out_read),
    .config_out_write(Tile_X01_Y0D_config_out_write),
    .config_read(Tile_X01_Y0C_config_out_read),
    .config_write(Tile_X01_Y0C_config_out_write),
    .hi(Tile_X01_Y0D_hi_unq1),
    .lo(Tile_X01_Y0D_lo_unq1),
    .read_config_data(Tile_X01_Y0D_read_config_data),
    .read_config_data_in(Tile_X01_Y0C_read_config_data),
    .reset(Tile_X01_Y0C_reset_out),
    .reset_out(Tile_X01_Y0D_reset_out),
    .stall(Tile_X01_Y0C_stall_out),
    .stall_out(Tile_X01_Y0D_stall_out),
    .tile_id(Tile_X01_Y0D_tile_id_in)
);
mantle_wire__typeBit9 Tile_X01_Y0D_hi (
    .in(Tile_X01_Y0D_hi_unq1),
    .out(Tile_X01_Y0D_hi_out)
);
mantle_wire__typeBit8 Tile_X01_Y0D_lo (
    .in(Tile_X01_Y0D_lo_unq1),
    .out(Tile_X01_Y0D_lo_out)
);
wire [15:0] Tile_X01_Y0D_tile_id_out;
assign Tile_X01_Y0D_tile_id_out = {Tile_X01_Y0D_lo_out[7],Tile_X01_Y0D_lo_out[7:6],Tile_X01_Y0D_lo_out[6:5],Tile_X01_Y0D_lo_out[5:4],Tile_X01_Y0D_hi_out[4],Tile_X01_Y0D_lo_out[3],Tile_X01_Y0D_lo_out[3:2],Tile_X01_Y0D_lo_out[2],Tile_X01_Y0D_hi_out[2:1],Tile_X01_Y0D_lo_out[0],Tile_X01_Y0D_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X01_Y0D_tile_id (
    .in(Tile_X01_Y0D_tile_id_in),
    .out(Tile_X01_Y0D_tile_id_out)
);
Tile_PE Tile_X01_Y0E (
    .SB_T0_EAST_SB_IN_B1(Tile_X02_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X02_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X01_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X01_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X01_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X00_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X00_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X01_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X02_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X02_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X01_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X01_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X01_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X00_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X00_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X01_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X02_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X02_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X01_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X01_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X01_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X00_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X00_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X01_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X02_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X02_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X01_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X01_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X01_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X01_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X01_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X01_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X01_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X00_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X00_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X01_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X02_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X02_Y0E_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X01_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X01_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X01_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X01_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X01_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X01_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X01_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X00_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X00_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X01_Y0E_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X01_Y0D_clk_out),
    .clk_out(Tile_X01_Y0E_clk_out),
    .clk_pass_through(Tile_X01_Y0D_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X01_Y0E_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X01_Y0E_clk_pass_through_out_right),
    .config_config_addr(Tile_X01_Y0D_config_out_config_addr),
    .config_config_data(Tile_X01_Y0D_config_out_config_data),
    .config_out_config_addr(Tile_X01_Y0E_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y0E_config_out_config_data),
    .config_out_read(Tile_X01_Y0E_config_out_read),
    .config_out_write(Tile_X01_Y0E_config_out_write),
    .config_read(Tile_X01_Y0D_config_out_read),
    .config_write(Tile_X01_Y0D_config_out_write),
    .hi(Tile_X01_Y0E_hi_unq1),
    .lo(Tile_X01_Y0E_lo_unq1),
    .read_config_data(Tile_X01_Y0E_read_config_data),
    .read_config_data_in(Tile_X01_Y0D_read_config_data),
    .reset(Tile_X01_Y0D_reset_out),
    .reset_out(Tile_X01_Y0E_reset_out),
    .stall(Tile_X01_Y0D_stall_out),
    .stall_out(Tile_X01_Y0E_stall_out),
    .tile_id(Tile_X01_Y0E_tile_id_in)
);
mantle_wire__typeBit9 Tile_X01_Y0E_hi (
    .in(Tile_X01_Y0E_hi_unq1),
    .out(Tile_X01_Y0E_hi_out)
);
mantle_wire__typeBit8 Tile_X01_Y0E_lo (
    .in(Tile_X01_Y0E_lo_unq1),
    .out(Tile_X01_Y0E_lo_out)
);
wire [15:0] Tile_X01_Y0E_tile_id_out;
assign Tile_X01_Y0E_tile_id_out = {Tile_X01_Y0E_lo_out[7],Tile_X01_Y0E_lo_out[7:6],Tile_X01_Y0E_lo_out[6:5],Tile_X01_Y0E_lo_out[5:4],Tile_X01_Y0E_hi_out[4],Tile_X01_Y0E_lo_out[3],Tile_X01_Y0E_lo_out[3:2],Tile_X01_Y0E_lo_out[2],Tile_X01_Y0E_hi_out[2:1],Tile_X01_Y0E_hi_out[1],Tile_X01_Y0E_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X01_Y0E_tile_id (
    .in(Tile_X01_Y0E_tile_id_in),
    .out(Tile_X01_Y0E_tile_id_out)
);
Tile_PE Tile_X01_Y0F (
    .SB_T0_EAST_SB_IN_B1(Tile_X02_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X02_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X01_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X01_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X01_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X01_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X01_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X00_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X00_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X01_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X02_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X02_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X01_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X01_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X01_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X01_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X01_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X00_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X00_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X01_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X02_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X02_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X01_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X01_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X01_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X01_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X01_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X00_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X00_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X01_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X02_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X02_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X01_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X01_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X01_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X01_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X01_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X01_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X01_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X00_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X00_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X01_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X02_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X02_Y0F_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X01_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X01_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X01_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X01_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X01_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X01_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X01_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X00_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X00_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X01_Y0F_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X01_Y0E_clk_out),
    .clk_out(Tile_X01_Y0F_clk_out),
    .clk_pass_through(Tile_X01_Y0E_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X01_Y0F_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X01_Y0F_clk_pass_through_out_right),
    .config_config_addr(Tile_X01_Y0E_config_out_config_addr),
    .config_config_data(Tile_X01_Y0E_config_out_config_data),
    .config_out_config_addr(Tile_X01_Y0F_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y0F_config_out_config_data),
    .config_out_read(Tile_X01_Y0F_config_out_read),
    .config_out_write(Tile_X01_Y0F_config_out_write),
    .config_read(Tile_X01_Y0E_config_out_read),
    .config_write(Tile_X01_Y0E_config_out_write),
    .hi(Tile_X01_Y0F_hi_unq1),
    .lo(Tile_X01_Y0F_lo_unq1),
    .read_config_data(Tile_X01_Y0F_read_config_data),
    .read_config_data_in(Tile_X01_Y0E_read_config_data),
    .reset(Tile_X01_Y0E_reset_out),
    .reset_out(Tile_X01_Y0F_reset_out),
    .stall(Tile_X01_Y0E_stall_out),
    .stall_out(Tile_X01_Y0F_stall_out),
    .tile_id(Tile_X01_Y0F_tile_id_in)
);
mantle_wire__typeBit9 Tile_X01_Y0F_hi (
    .in(Tile_X01_Y0F_hi_unq1),
    .out(Tile_X01_Y0F_hi_out)
);
mantle_wire__typeBit8 Tile_X01_Y0F_lo (
    .in(Tile_X01_Y0F_lo_unq1),
    .out(Tile_X01_Y0F_lo_out)
);
wire [15:0] Tile_X01_Y0F_tile_id_out;
assign Tile_X01_Y0F_tile_id_out = {Tile_X01_Y0F_lo_out[7],Tile_X01_Y0F_lo_out[7:6],Tile_X01_Y0F_lo_out[6:5],Tile_X01_Y0F_lo_out[5:4],Tile_X01_Y0F_hi_out[4],Tile_X01_Y0F_lo_out[3],Tile_X01_Y0F_lo_out[3:2],Tile_X01_Y0F_lo_out[2],Tile_X01_Y0F_hi_out[2:1],Tile_X01_Y0F_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X01_Y0F_tile_id (
    .in(Tile_X01_Y0F_tile_id_in),
    .out(Tile_X01_Y0F_tile_id_out)
);
Tile_PE Tile_X01_Y10 (
    .SB_T0_EAST_SB_IN_B1(Tile_X02_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X02_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X01_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X01_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X01_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X01_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X01_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X01_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T0_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X01_Y10_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X01_Y10_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X00_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X00_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X01_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X01_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X02_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X02_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X01_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X01_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X01_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X01_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X01_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X01_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T1_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X01_Y10_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X01_Y10_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X00_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X00_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X01_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X01_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X02_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X02_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X01_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X01_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X01_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X01_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X01_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X01_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T2_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X01_Y10_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X01_Y10_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X00_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X00_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X01_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X01_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X02_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X02_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X01_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X01_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X01_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X01_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X01_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X01_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T3_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X01_Y10_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X01_Y10_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X00_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X00_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X01_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X01_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X02_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X02_Y10_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X01_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X01_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X01_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X01_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X01_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X01_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T4_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X01_Y10_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X01_Y10_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X00_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X00_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X01_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X01_Y10_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X01_Y0F_clk_out),
    .clk_out(Tile_X01_Y10_clk_out),
    .clk_pass_through(Tile_X01_Y0F_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X01_Y10_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X01_Y10_clk_pass_through_out_right),
    .config_config_addr(Tile_X01_Y0F_config_out_config_addr),
    .config_config_data(Tile_X01_Y0F_config_out_config_data),
    .config_out_config_addr(Tile_X01_Y10_config_out_config_addr),
    .config_out_config_data(Tile_X01_Y10_config_out_config_data),
    .config_out_read(Tile_X01_Y10_config_out_read),
    .config_out_write(Tile_X01_Y10_config_out_write),
    .config_read(Tile_X01_Y0F_config_out_read),
    .config_write(Tile_X01_Y0F_config_out_write),
    .hi(Tile_X01_Y10_hi),
    .lo(Tile_X01_Y10_lo_unq1),
    .read_config_data(Tile_X01_Y10_read_config_data),
    .read_config_data_in(Tile_X01_Y0F_read_config_data),
    .reset(Tile_X01_Y0F_reset_out),
    .reset_out(Tile_X01_Y10_reset_out),
    .stall(Tile_X01_Y0F_stall_out),
    .stall_out(Tile_X01_Y10_stall_out),
    .tile_id(Tile_X01_Y10_tile_id_in)
);
mantle_wire__typeBit8 Tile_X01_Y10_lo (
    .in(Tile_X01_Y10_lo_unq1),
    .out(Tile_X01_Y10_lo_out)
);
wire [15:0] Tile_X01_Y10_tile_id_out;
assign Tile_X01_Y10_tile_id_out = {Tile_X01_Y10_lo_out[7],Tile_X01_Y10_lo_out[7:6],Tile_X01_Y10_lo_out[6:5],Tile_X01_Y10_lo_out[5:4],Tile_X01_Y10_hi[4],Tile_X01_Y10_lo_out[3],Tile_X01_Y10_lo_out[3:2],Tile_X01_Y10_hi[2],Tile_X01_Y10_lo_out[1],Tile_X01_Y10_lo_out[1:0],Tile_X01_Y10_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X01_Y10_tile_id (
    .in(Tile_X01_Y10_tile_id_in),
    .out(Tile_X01_Y10_tile_id_out)
);
wire [15:0] Tile_X02_Y00_tile_id;
assign Tile_X02_Y00_tile_id = {Tile_X02_Y00_lo[7],Tile_X02_Y00_lo[7:6],Tile_X02_Y00_lo[6:5],Tile_X02_Y00_lo[5],Tile_X02_Y00_hi[5],Tile_X02_Y00_lo[4:3],Tile_X02_Y00_lo[3:2],Tile_X02_Y00_lo[2:1],Tile_X02_Y00_lo[1:0],Tile_X02_Y00_lo[0]};
Tile_io_core Tile_X02_Y00 (
    .tile_id(Tile_X02_Y00_tile_id),
    .glb2io_1(glb2io_1_X02_Y00),
    .f2io_1(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B1),
    .io2glb_1(Tile_X02_Y00_io2glb_1),
    .io2f_1(Tile_X02_Y00_io2f_1),
    .glb2io_16(glb2io_16_X02_Y00),
    .f2io_16(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B16),
    .io2glb_16(Tile_X02_Y00_io2glb_16),
    .io2f_16(Tile_X02_Y00_io2f_16),
    .hi(Tile_X02_Y00_hi),
    .lo(Tile_X02_Y00_lo)
);
Tile_PE Tile_X02_Y01 (
    .SB_T0_EAST_SB_IN_B1(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X02_Y00_io2f_1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X02_Y00_io2f_16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y01_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X01_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X02_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X02_Y00_io2f_1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X02_Y00_io2f_16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y01_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X01_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X02_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X02_Y00_io2f_1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X02_Y00_io2f_16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y01_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X01_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X02_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X03_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X03_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X02_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X02_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X02_Y00_io2f_1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X02_Y00_io2f_16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y01_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X02_Y01_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X01_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X01_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X02_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X02_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X03_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X03_Y01_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X02_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X02_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X02_Y00_io2f_1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X02_Y00_io2f_16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y01_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X02_Y01_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X01_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X01_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X02_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X02_Y01_SB_T4_WEST_SB_OUT_B16),
    .clk(clk),
    .clk_out(Tile_X02_Y01_clk_out),
    .clk_pass_through(clk),
    .clk_pass_through_out_bot(Tile_X02_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X02_Y01_clk_pass_through_out_right),
    .config_config_addr(config_2_config_addr),
    .config_config_data(config_2_config_data),
    .config_out_config_addr(Tile_X02_Y01_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y01_config_out_config_data),
    .config_out_read(Tile_X02_Y01_config_out_read),
    .config_out_write(Tile_X02_Y01_config_out_write),
    .config_read(config_2_read),
    .config_write(config_2_write),
    .hi(Tile_X02_Y01_hi),
    .lo(Tile_X02_Y01_lo_unq1),
    .read_config_data(Tile_X02_Y01_read_config_data),
    .read_config_data_in(const_0_32_out),
    .reset(reset),
    .reset_out(Tile_X02_Y01_reset_out),
    .stall(stall[2]),
    .stall_out(Tile_X02_Y01_stall_out),
    .tile_id(Tile_X02_Y01_tile_id_in)
);
mantle_wire__typeBit8 Tile_X02_Y01_lo (
    .in(Tile_X02_Y01_lo_unq1),
    .out(Tile_X02_Y01_lo_out)
);
wire [15:0] Tile_X02_Y01_tile_id_out;
assign Tile_X02_Y01_tile_id_out = {Tile_X02_Y01_lo_out[7],Tile_X02_Y01_lo_out[7:6],Tile_X02_Y01_lo_out[6:5],Tile_X02_Y01_lo_out[5],Tile_X02_Y01_hi[5],Tile_X02_Y01_lo_out[4:3],Tile_X02_Y01_lo_out[3:2],Tile_X02_Y01_lo_out[2:1],Tile_X02_Y01_lo_out[1:0],Tile_X02_Y01_hi[0]};
mantle_wire__typeBitIn16 Tile_X02_Y01_tile_id (
    .in(Tile_X02_Y01_tile_id_in),
    .out(Tile_X02_Y01_tile_id_out)
);
Tile_PE Tile_X02_Y02 (
    .SB_T0_EAST_SB_IN_B1(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X02_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X01_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X02_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X02_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X01_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X02_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X02_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X01_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X02_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X03_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X03_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X02_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X02_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X02_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X02_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X01_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X01_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X02_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X02_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X03_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X03_Y02_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X02_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X02_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X02_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X02_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X01_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X01_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X02_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X02_Y02_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y01_clk_out),
    .clk_out(Tile_X02_Y02_clk_out),
    .clk_pass_through(Tile_X02_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X02_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X02_Y02_clk_pass_through_out_right),
    .config_config_addr(Tile_X02_Y01_config_out_config_addr),
    .config_config_data(Tile_X02_Y01_config_out_config_data),
    .config_out_config_addr(Tile_X02_Y02_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y02_config_out_config_data),
    .config_out_read(Tile_X02_Y02_config_out_read),
    .config_out_write(Tile_X02_Y02_config_out_write),
    .config_read(Tile_X02_Y01_config_out_read),
    .config_write(Tile_X02_Y01_config_out_write),
    .hi(Tile_X02_Y02_hi),
    .lo(Tile_X02_Y02_lo_unq1),
    .read_config_data(Tile_X02_Y02_read_config_data),
    .read_config_data_in(Tile_X02_Y01_read_config_data),
    .reset(Tile_X02_Y01_reset_out),
    .reset_out(Tile_X02_Y02_reset_out),
    .stall(Tile_X02_Y01_stall_out),
    .stall_out(Tile_X02_Y02_stall_out),
    .tile_id(Tile_X02_Y02_tile_id_in)
);
mantle_wire__typeBit8 Tile_X02_Y02_lo (
    .in(Tile_X02_Y02_lo_unq1),
    .out(Tile_X02_Y02_lo_out)
);
wire [15:0] Tile_X02_Y02_tile_id_out;
assign Tile_X02_Y02_tile_id_out = {Tile_X02_Y02_lo_out[7],Tile_X02_Y02_lo_out[7:6],Tile_X02_Y02_lo_out[6:5],Tile_X02_Y02_lo_out[5],Tile_X02_Y02_hi[5],Tile_X02_Y02_lo_out[4:3],Tile_X02_Y02_lo_out[3:2],Tile_X02_Y02_lo_out[2:1],Tile_X02_Y02_lo_out[1],Tile_X02_Y02_hi[1],Tile_X02_Y02_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X02_Y02_tile_id (
    .in(Tile_X02_Y02_tile_id_in),
    .out(Tile_X02_Y02_tile_id_out)
);
Tile_PE Tile_X02_Y03 (
    .SB_T0_EAST_SB_IN_B1(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X02_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X01_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X02_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X02_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X01_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X02_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X02_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X01_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X02_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X03_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X03_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X02_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X02_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X02_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X02_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X01_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X01_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X02_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X02_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X03_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X03_Y03_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X02_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X02_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X02_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X02_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X01_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X01_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X02_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X02_Y03_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y02_clk_out),
    .clk_out(Tile_X02_Y03_clk_out),
    .clk_pass_through(Tile_X02_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X02_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X02_Y03_clk_pass_through_out_right),
    .config_config_addr(Tile_X02_Y02_config_out_config_addr),
    .config_config_data(Tile_X02_Y02_config_out_config_data),
    .config_out_config_addr(Tile_X02_Y03_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y03_config_out_config_data),
    .config_out_read(Tile_X02_Y03_config_out_read),
    .config_out_write(Tile_X02_Y03_config_out_write),
    .config_read(Tile_X02_Y02_config_out_read),
    .config_write(Tile_X02_Y02_config_out_write),
    .hi(Tile_X02_Y03_hi_unq1),
    .lo(Tile_X02_Y03_lo_unq1),
    .read_config_data(Tile_X02_Y03_read_config_data),
    .read_config_data_in(Tile_X02_Y02_read_config_data),
    .reset(Tile_X02_Y02_reset_out),
    .reset_out(Tile_X02_Y03_reset_out),
    .stall(Tile_X02_Y02_stall_out),
    .stall_out(Tile_X02_Y03_stall_out),
    .tile_id(Tile_X02_Y03_tile_id_in)
);
mantle_wire__typeBit9 Tile_X02_Y03_hi (
    .in(Tile_X02_Y03_hi_unq1),
    .out(Tile_X02_Y03_hi_out)
);
mantle_wire__typeBit8 Tile_X02_Y03_lo (
    .in(Tile_X02_Y03_lo_unq1),
    .out(Tile_X02_Y03_lo_out)
);
wire [15:0] Tile_X02_Y03_tile_id_out;
assign Tile_X02_Y03_tile_id_out = {Tile_X02_Y03_lo_out[7],Tile_X02_Y03_lo_out[7:6],Tile_X02_Y03_lo_out[6:5],Tile_X02_Y03_lo_out[5],Tile_X02_Y03_hi_out[5],Tile_X02_Y03_lo_out[4:3],Tile_X02_Y03_lo_out[3:2],Tile_X02_Y03_lo_out[2:1],Tile_X02_Y03_lo_out[1],Tile_X02_Y03_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X02_Y03_tile_id (
    .in(Tile_X02_Y03_tile_id_in),
    .out(Tile_X02_Y03_tile_id_out)
);
Tile_PE Tile_X02_Y04 (
    .SB_T0_EAST_SB_IN_B1(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X02_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X01_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X02_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X02_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X01_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X02_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X02_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X01_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X02_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X03_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X03_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X02_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X02_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X02_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X02_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X02_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X02_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X01_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X01_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X02_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X02_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X03_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X03_Y04_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X02_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X02_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X02_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X02_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X02_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X02_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X01_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X01_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X02_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X02_Y04_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y03_clk_out),
    .clk_out(Tile_X02_Y04_clk_out),
    .clk_pass_through(Tile_X02_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X02_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X02_Y04_clk_pass_through_out_right),
    .config_config_addr(Tile_X02_Y03_config_out_config_addr),
    .config_config_data(Tile_X02_Y03_config_out_config_data),
    .config_out_config_addr(Tile_X02_Y04_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y04_config_out_config_data),
    .config_out_read(Tile_X02_Y04_config_out_read),
    .config_out_write(Tile_X02_Y04_config_out_write),
    .config_read(Tile_X02_Y03_config_out_read),
    .config_write(Tile_X02_Y03_config_out_write),
    .hi(Tile_X02_Y04_hi),
    .lo(Tile_X02_Y04_lo_unq1),
    .read_config_data(Tile_X02_Y04_read_config_data),
    .read_config_data_in(Tile_X02_Y03_read_config_data),
    .reset(Tile_X02_Y03_reset_out),
    .reset_out(Tile_X02_Y04_reset_out),
    .stall(Tile_X02_Y03_stall_out),
    .stall_out(Tile_X02_Y04_stall_out),
    .tile_id(Tile_X02_Y04_tile_id_in)
);
mantle_wire__typeBit8 Tile_X02_Y04_lo (
    .in(Tile_X02_Y04_lo_unq1),
    .out(Tile_X02_Y04_lo_out)
);
wire [15:0] Tile_X02_Y04_tile_id_out;
assign Tile_X02_Y04_tile_id_out = {Tile_X02_Y04_lo_out[7],Tile_X02_Y04_lo_out[7:6],Tile_X02_Y04_lo_out[6:5],Tile_X02_Y04_lo_out[5],Tile_X02_Y04_hi[5],Tile_X02_Y04_lo_out[4:3],Tile_X02_Y04_lo_out[3:2],Tile_X02_Y04_lo_out[2:1],Tile_X02_Y04_hi[1],Tile_X02_Y04_lo_out[0],Tile_X02_Y04_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X02_Y04_tile_id (
    .in(Tile_X02_Y04_tile_id_in),
    .out(Tile_X02_Y04_tile_id_out)
);
Tile_PE Tile_X02_Y05 (
    .SB_T0_EAST_SB_IN_B1(Tile_X03_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X03_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X02_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X02_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X02_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X01_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X01_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X02_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X02_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X03_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X03_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X02_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X02_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X02_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X01_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X01_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X02_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X02_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X03_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X03_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X02_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X02_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X02_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X01_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X01_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X02_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X02_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X03_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X03_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X02_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X02_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X02_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X02_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X02_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X02_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X02_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X01_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X01_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X02_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X02_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X03_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X03_Y05_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X02_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X02_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X02_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X02_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X02_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X02_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X02_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X01_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X01_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X02_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X02_Y05_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y04_clk_out),
    .clk_out(Tile_X02_Y05_clk_out),
    .clk_pass_through(Tile_X02_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X02_Y05_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X02_Y05_clk_pass_through_out_right),
    .config_config_addr(Tile_X02_Y04_config_out_config_addr),
    .config_config_data(Tile_X02_Y04_config_out_config_data),
    .config_out_config_addr(Tile_X02_Y05_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y05_config_out_config_data),
    .config_out_read(Tile_X02_Y05_config_out_read),
    .config_out_write(Tile_X02_Y05_config_out_write),
    .config_read(Tile_X02_Y04_config_out_read),
    .config_write(Tile_X02_Y04_config_out_write),
    .hi(Tile_X02_Y05_hi),
    .lo(Tile_X02_Y05_lo_unq1),
    .read_config_data(Tile_X02_Y05_read_config_data),
    .read_config_data_in(Tile_X02_Y04_read_config_data),
    .reset(Tile_X02_Y04_reset_out),
    .reset_out(Tile_X02_Y05_reset_out),
    .stall(Tile_X02_Y04_stall_out),
    .stall_out(Tile_X02_Y05_stall_out),
    .tile_id(Tile_X02_Y05_tile_id_in)
);
mantle_wire__typeBit8 Tile_X02_Y05_lo (
    .in(Tile_X02_Y05_lo_unq1),
    .out(Tile_X02_Y05_lo_out)
);
wire [15:0] Tile_X02_Y05_tile_id_out;
assign Tile_X02_Y05_tile_id_out = {Tile_X02_Y05_lo_out[7],Tile_X02_Y05_lo_out[7:6],Tile_X02_Y05_lo_out[6:5],Tile_X02_Y05_lo_out[5],Tile_X02_Y05_hi[5],Tile_X02_Y05_lo_out[4:3],Tile_X02_Y05_lo_out[3:2],Tile_X02_Y05_lo_out[2:1],Tile_X02_Y05_hi[1],Tile_X02_Y05_lo_out[0],Tile_X02_Y05_hi[0]};
mantle_wire__typeBitIn16 Tile_X02_Y05_tile_id (
    .in(Tile_X02_Y05_tile_id_in),
    .out(Tile_X02_Y05_tile_id_out)
);
Tile_PE Tile_X02_Y06 (
    .SB_T0_EAST_SB_IN_B1(Tile_X03_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X03_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X02_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X02_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X02_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X02_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X01_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X01_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X02_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X02_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X03_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X03_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X02_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X02_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X02_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X02_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X01_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X01_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X02_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X02_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X03_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X03_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X02_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X02_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X02_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X02_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X01_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X01_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X02_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X02_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X03_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X03_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X02_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X02_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X02_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X02_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X02_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X02_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X02_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X02_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X01_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X01_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X02_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X02_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X03_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X03_Y06_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X02_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X02_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X02_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X02_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X02_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X02_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X02_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X02_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X01_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X01_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X02_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X02_Y06_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y05_clk_out),
    .clk_out(Tile_X02_Y06_clk_out),
    .clk_pass_through(Tile_X02_Y05_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X02_Y06_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X02_Y06_clk_pass_through_out_right),
    .config_config_addr(Tile_X02_Y05_config_out_config_addr),
    .config_config_data(Tile_X02_Y05_config_out_config_data),
    .config_out_config_addr(Tile_X02_Y06_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y06_config_out_config_data),
    .config_out_read(Tile_X02_Y06_config_out_read),
    .config_out_write(Tile_X02_Y06_config_out_write),
    .config_read(Tile_X02_Y05_config_out_read),
    .config_write(Tile_X02_Y05_config_out_write),
    .hi(Tile_X02_Y06_hi),
    .lo(Tile_X02_Y06_lo_unq1),
    .read_config_data(Tile_X02_Y06_read_config_data),
    .read_config_data_in(Tile_X02_Y05_read_config_data),
    .reset(Tile_X02_Y05_reset_out),
    .reset_out(Tile_X02_Y06_reset_out),
    .stall(Tile_X02_Y05_stall_out),
    .stall_out(Tile_X02_Y06_stall_out),
    .tile_id(Tile_X02_Y06_tile_id_in)
);
mantle_wire__typeBit8 Tile_X02_Y06_lo (
    .in(Tile_X02_Y06_lo_unq1),
    .out(Tile_X02_Y06_lo_out)
);
wire [15:0] Tile_X02_Y06_tile_id_out;
assign Tile_X02_Y06_tile_id_out = {Tile_X02_Y06_lo_out[7],Tile_X02_Y06_lo_out[7:6],Tile_X02_Y06_lo_out[6:5],Tile_X02_Y06_lo_out[5],Tile_X02_Y06_hi[5],Tile_X02_Y06_lo_out[4:3],Tile_X02_Y06_lo_out[3:2],Tile_X02_Y06_lo_out[2:1],Tile_X02_Y06_hi[1],Tile_X02_Y06_hi[1],Tile_X02_Y06_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X02_Y06_tile_id (
    .in(Tile_X02_Y06_tile_id_in),
    .out(Tile_X02_Y06_tile_id_out)
);
Tile_PE Tile_X02_Y07 (
    .SB_T0_EAST_SB_IN_B1(Tile_X03_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X03_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X02_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X02_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X02_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X02_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X01_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X01_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X02_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X02_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X03_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X03_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X02_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X02_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X02_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X02_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X01_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X01_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X02_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X02_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X03_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X03_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X02_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X02_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X02_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X02_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X01_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X01_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X02_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X02_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X03_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X03_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X02_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X02_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X02_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X02_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X02_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X02_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X02_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X02_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X01_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X01_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X02_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X02_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X03_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X03_Y07_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X02_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X02_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X02_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X02_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X02_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X02_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X02_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X02_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X01_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X01_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X02_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X02_Y07_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y06_clk_out),
    .clk_out(Tile_X02_Y07_clk_out),
    .clk_pass_through(Tile_X02_Y06_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X02_Y07_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X02_Y07_clk_pass_through_out_right),
    .config_config_addr(Tile_X02_Y06_config_out_config_addr),
    .config_config_data(Tile_X02_Y06_config_out_config_data),
    .config_out_config_addr(Tile_X02_Y07_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y07_config_out_config_data),
    .config_out_read(Tile_X02_Y07_config_out_read),
    .config_out_write(Tile_X02_Y07_config_out_write),
    .config_read(Tile_X02_Y06_config_out_read),
    .config_write(Tile_X02_Y06_config_out_write),
    .hi(Tile_X02_Y07_hi_unq1),
    .lo(Tile_X02_Y07_lo_unq1),
    .read_config_data(Tile_X02_Y07_read_config_data),
    .read_config_data_in(Tile_X02_Y06_read_config_data),
    .reset(Tile_X02_Y06_reset_out),
    .reset_out(Tile_X02_Y07_reset_out),
    .stall(Tile_X02_Y06_stall_out),
    .stall_out(Tile_X02_Y07_stall_out),
    .tile_id(Tile_X02_Y07_tile_id_in)
);
mantle_wire__typeBit9 Tile_X02_Y07_hi (
    .in(Tile_X02_Y07_hi_unq1),
    .out(Tile_X02_Y07_hi_out)
);
mantle_wire__typeBit8 Tile_X02_Y07_lo (
    .in(Tile_X02_Y07_lo_unq1),
    .out(Tile_X02_Y07_lo_out)
);
wire [15:0] Tile_X02_Y07_tile_id_out;
assign Tile_X02_Y07_tile_id_out = {Tile_X02_Y07_lo_out[7],Tile_X02_Y07_lo_out[7:6],Tile_X02_Y07_lo_out[6:5],Tile_X02_Y07_lo_out[5],Tile_X02_Y07_hi_out[5],Tile_X02_Y07_lo_out[4:3],Tile_X02_Y07_lo_out[3:2],Tile_X02_Y07_lo_out[2:1],Tile_X02_Y07_hi_out[1],Tile_X02_Y07_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X02_Y07_tile_id (
    .in(Tile_X02_Y07_tile_id_in),
    .out(Tile_X02_Y07_tile_id_out)
);
Tile_PE Tile_X02_Y08 (
    .SB_T0_EAST_SB_IN_B1(Tile_X03_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X03_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X02_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X02_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X02_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X02_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X01_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X01_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X02_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X02_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X03_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X03_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X02_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X02_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X02_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X02_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X01_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X01_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X02_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X02_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X03_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X03_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X02_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X02_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X02_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X02_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X01_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X01_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X02_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X02_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X03_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X03_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X02_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X02_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X02_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X02_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X02_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X02_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X02_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X02_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X01_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X01_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X02_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X02_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X03_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X03_Y08_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X02_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X02_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X02_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X02_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X02_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X02_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X02_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X02_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X01_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X01_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X02_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X02_Y08_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y07_clk_out),
    .clk_out(Tile_X02_Y08_clk_out),
    .clk_pass_through(Tile_X02_Y07_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X02_Y08_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X02_Y08_clk_pass_through_out_right),
    .config_config_addr(Tile_X02_Y07_config_out_config_addr),
    .config_config_data(Tile_X02_Y07_config_out_config_data),
    .config_out_config_addr(Tile_X02_Y08_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y08_config_out_config_data),
    .config_out_read(Tile_X02_Y08_config_out_read),
    .config_out_write(Tile_X02_Y08_config_out_write),
    .config_read(Tile_X02_Y07_config_out_read),
    .config_write(Tile_X02_Y07_config_out_write),
    .hi(Tile_X02_Y08_hi),
    .lo(Tile_X02_Y08_lo_unq1),
    .read_config_data(Tile_X02_Y08_read_config_data),
    .read_config_data_in(Tile_X02_Y07_read_config_data),
    .reset(Tile_X02_Y07_reset_out),
    .reset_out(Tile_X02_Y08_reset_out),
    .stall(Tile_X02_Y07_stall_out),
    .stall_out(Tile_X02_Y08_stall_out),
    .tile_id(Tile_X02_Y08_tile_id_in)
);
mantle_wire__typeBit8 Tile_X02_Y08_lo (
    .in(Tile_X02_Y08_lo_unq1),
    .out(Tile_X02_Y08_lo_out)
);
wire [15:0] Tile_X02_Y08_tile_id_out;
assign Tile_X02_Y08_tile_id_out = {Tile_X02_Y08_lo_out[7],Tile_X02_Y08_lo_out[7:6],Tile_X02_Y08_lo_out[6:5],Tile_X02_Y08_lo_out[5],Tile_X02_Y08_hi[5],Tile_X02_Y08_lo_out[4:3],Tile_X02_Y08_lo_out[3:2],Tile_X02_Y08_lo_out[2],Tile_X02_Y08_hi[2],Tile_X02_Y08_lo_out[1:0],Tile_X02_Y08_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X02_Y08_tile_id (
    .in(Tile_X02_Y08_tile_id_in),
    .out(Tile_X02_Y08_tile_id_out)
);
Tile_PE Tile_X02_Y09 (
    .SB_T0_EAST_SB_IN_B1(Tile_X03_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X03_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X02_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X02_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X02_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X02_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X01_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X01_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X02_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X02_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X03_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X03_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X02_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X02_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X02_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X02_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X01_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X01_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X02_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X02_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X03_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X03_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X02_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X02_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X02_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X02_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X01_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X01_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X02_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X02_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X03_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X03_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X02_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X02_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X02_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X02_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X02_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X02_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X02_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X02_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X01_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X01_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X02_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X02_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X03_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X03_Y09_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X02_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X02_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X02_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X02_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X02_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X02_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X02_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X02_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X01_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X01_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X02_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X02_Y09_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y08_clk_out),
    .clk_out(Tile_X02_Y09_clk_out),
    .clk_pass_through(Tile_X02_Y08_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X02_Y09_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X02_Y09_clk_pass_through_out_right),
    .config_config_addr(ConfigPipeStage_inst2_config_out_config_addr),
    .config_config_data(ConfigPipeStage_inst2_config_out_config_data),
    .config_out_config_addr(Tile_X02_Y09_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y09_config_out_config_data),
    .config_out_read(Tile_X02_Y09_config_out_read),
    .config_out_write(Tile_X02_Y09_config_out_write),
    .config_read(ConfigPipeStage_inst2_config_out_read),
    .config_write(ConfigPipeStage_inst2_config_out_write),
    .hi(Tile_X02_Y09_hi),
    .lo(Tile_X02_Y09_lo_unq1),
    .read_config_data(Tile_X02_Y09_read_config_data),
    .read_config_data_in(Tile_X02_Y08_read_config_data),
    .reset(Tile_X02_Y08_reset_out),
    .reset_out(Tile_X02_Y09_reset_out),
    .stall(Tile_X02_Y08_stall_out),
    .stall_out(Tile_X02_Y09_stall_out),
    .tile_id(Tile_X02_Y09_tile_id_in)
);
mantle_wire__typeBit8 Tile_X02_Y09_lo (
    .in(Tile_X02_Y09_lo_unq1),
    .out(Tile_X02_Y09_lo_out)
);
wire [15:0] Tile_X02_Y09_tile_id_out;
assign Tile_X02_Y09_tile_id_out = {Tile_X02_Y09_lo_out[7],Tile_X02_Y09_lo_out[7:6],Tile_X02_Y09_lo_out[6:5],Tile_X02_Y09_lo_out[5],Tile_X02_Y09_hi[5],Tile_X02_Y09_lo_out[4:3],Tile_X02_Y09_lo_out[3:2],Tile_X02_Y09_lo_out[2],Tile_X02_Y09_hi[2],Tile_X02_Y09_lo_out[1:0],Tile_X02_Y09_hi[0]};
mantle_wire__typeBitIn16 Tile_X02_Y09_tile_id (
    .in(Tile_X02_Y09_tile_id_in),
    .out(Tile_X02_Y09_tile_id_out)
);
Tile_PE Tile_X02_Y0A (
    .SB_T0_EAST_SB_IN_B1(Tile_X03_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X03_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X02_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X02_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X02_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X02_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X01_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X01_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X02_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X02_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X03_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X03_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X02_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X02_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X02_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X02_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X01_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X01_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X02_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X02_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X03_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X03_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X02_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X02_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X02_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X02_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X01_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X01_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X02_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X02_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X03_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X03_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X02_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X02_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X02_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X02_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X02_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X02_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X02_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X02_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X01_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X01_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X02_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X02_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X03_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X03_Y0A_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X02_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X02_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X02_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X02_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X02_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X02_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X02_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X02_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X01_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X01_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X02_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X02_Y0A_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y09_clk_out),
    .clk_out(Tile_X02_Y0A_clk_out),
    .clk_pass_through(Tile_X02_Y09_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X02_Y0A_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X02_Y0A_clk_pass_through_out_right),
    .config_config_addr(Tile_X02_Y09_config_out_config_addr),
    .config_config_data(Tile_X02_Y09_config_out_config_data),
    .config_out_config_addr(Tile_X02_Y0A_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y0A_config_out_config_data),
    .config_out_read(Tile_X02_Y0A_config_out_read),
    .config_out_write(Tile_X02_Y0A_config_out_write),
    .config_read(Tile_X02_Y09_config_out_read),
    .config_write(Tile_X02_Y09_config_out_write),
    .hi(Tile_X02_Y0A_hi),
    .lo(Tile_X02_Y0A_lo_unq1),
    .read_config_data(Tile_X02_Y0A_read_config_data),
    .read_config_data_in(Tile_X02_Y09_read_config_data),
    .reset(Tile_X02_Y09_reset_out),
    .reset_out(Tile_X02_Y0A_reset_out),
    .stall(Tile_X02_Y09_stall_out),
    .stall_out(Tile_X02_Y0A_stall_out),
    .tile_id(Tile_X02_Y0A_tile_id_in)
);
mantle_wire__typeBit8 Tile_X02_Y0A_lo (
    .in(Tile_X02_Y0A_lo_unq1),
    .out(Tile_X02_Y0A_lo_out)
);
wire [15:0] Tile_X02_Y0A_tile_id_out;
assign Tile_X02_Y0A_tile_id_out = {Tile_X02_Y0A_lo_out[7],Tile_X02_Y0A_lo_out[7:6],Tile_X02_Y0A_lo_out[6:5],Tile_X02_Y0A_lo_out[5],Tile_X02_Y0A_hi[5],Tile_X02_Y0A_lo_out[4:3],Tile_X02_Y0A_lo_out[3:2],Tile_X02_Y0A_lo_out[2],Tile_X02_Y0A_hi[2],Tile_X02_Y0A_lo_out[1],Tile_X02_Y0A_hi[1],Tile_X02_Y0A_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X02_Y0A_tile_id (
    .in(Tile_X02_Y0A_tile_id_in),
    .out(Tile_X02_Y0A_tile_id_out)
);
Tile_PE Tile_X02_Y0B (
    .SB_T0_EAST_SB_IN_B1(Tile_X03_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X03_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X02_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X02_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X02_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X02_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X01_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X01_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X02_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X02_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X03_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X03_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X02_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X02_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X02_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X02_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X01_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X01_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X02_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X02_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X03_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X03_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X02_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X02_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X02_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X02_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X01_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X01_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X02_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X02_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X03_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X03_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X02_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X02_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X02_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X02_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X02_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X02_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X02_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X02_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X01_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X01_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X02_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X02_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X03_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X03_Y0B_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X02_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X02_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X02_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X02_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X02_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X02_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X02_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X02_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X01_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X01_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X02_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X02_Y0B_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y0A_clk_out),
    .clk_out(Tile_X02_Y0B_clk_out),
    .clk_pass_through(Tile_X02_Y0A_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X02_Y0B_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X02_Y0B_clk_pass_through_out_right),
    .config_config_addr(Tile_X02_Y0A_config_out_config_addr),
    .config_config_data(Tile_X02_Y0A_config_out_config_data),
    .config_out_config_addr(Tile_X02_Y0B_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y0B_config_out_config_data),
    .config_out_read(Tile_X02_Y0B_config_out_read),
    .config_out_write(Tile_X02_Y0B_config_out_write),
    .config_read(Tile_X02_Y0A_config_out_read),
    .config_write(Tile_X02_Y0A_config_out_write),
    .hi(Tile_X02_Y0B_hi_unq1),
    .lo(Tile_X02_Y0B_lo_unq1),
    .read_config_data(Tile_X02_Y0B_read_config_data),
    .read_config_data_in(Tile_X02_Y0A_read_config_data),
    .reset(Tile_X02_Y0A_reset_out),
    .reset_out(Tile_X02_Y0B_reset_out),
    .stall(Tile_X02_Y0A_stall_out),
    .stall_out(Tile_X02_Y0B_stall_out),
    .tile_id(Tile_X02_Y0B_tile_id_in)
);
mantle_wire__typeBit9 Tile_X02_Y0B_hi (
    .in(Tile_X02_Y0B_hi_unq1),
    .out(Tile_X02_Y0B_hi_out)
);
mantle_wire__typeBit8 Tile_X02_Y0B_lo (
    .in(Tile_X02_Y0B_lo_unq1),
    .out(Tile_X02_Y0B_lo_out)
);
wire [15:0] Tile_X02_Y0B_tile_id_out;
assign Tile_X02_Y0B_tile_id_out = {Tile_X02_Y0B_lo_out[7],Tile_X02_Y0B_lo_out[7:6],Tile_X02_Y0B_lo_out[6:5],Tile_X02_Y0B_lo_out[5],Tile_X02_Y0B_hi_out[5],Tile_X02_Y0B_lo_out[4:3],Tile_X02_Y0B_lo_out[3:2],Tile_X02_Y0B_lo_out[2],Tile_X02_Y0B_hi_out[2],Tile_X02_Y0B_lo_out[1],Tile_X02_Y0B_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X02_Y0B_tile_id (
    .in(Tile_X02_Y0B_tile_id_in),
    .out(Tile_X02_Y0B_tile_id_out)
);
Tile_PE Tile_X02_Y0C (
    .SB_T0_EAST_SB_IN_B1(Tile_X03_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X03_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X02_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X02_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X02_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X02_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X01_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X01_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X02_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X02_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X03_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X03_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X02_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X02_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X02_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X02_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X01_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X01_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X02_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X02_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X03_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X03_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X02_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X02_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X02_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X02_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X01_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X01_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X02_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X02_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X03_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X03_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X02_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X02_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X02_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X02_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X02_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X02_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X02_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X02_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X01_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X01_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X02_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X02_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X03_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X03_Y0C_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X02_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X02_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X02_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X02_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X02_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X02_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X02_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X02_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X01_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X01_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X02_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X02_Y0C_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y0B_clk_out),
    .clk_out(Tile_X02_Y0C_clk_out),
    .clk_pass_through(Tile_X02_Y0B_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X02_Y0C_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X02_Y0C_clk_pass_through_out_right),
    .config_config_addr(Tile_X02_Y0B_config_out_config_addr),
    .config_config_data(Tile_X02_Y0B_config_out_config_data),
    .config_out_config_addr(Tile_X02_Y0C_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y0C_config_out_config_data),
    .config_out_read(Tile_X02_Y0C_config_out_read),
    .config_out_write(Tile_X02_Y0C_config_out_write),
    .config_read(Tile_X02_Y0B_config_out_read),
    .config_write(Tile_X02_Y0B_config_out_write),
    .hi(Tile_X02_Y0C_hi_unq1),
    .lo(Tile_X02_Y0C_lo_unq1),
    .read_config_data(Tile_X02_Y0C_read_config_data),
    .read_config_data_in(Tile_X02_Y0B_read_config_data),
    .reset(Tile_X02_Y0B_reset_out),
    .reset_out(Tile_X02_Y0C_reset_out),
    .stall(Tile_X02_Y0B_stall_out),
    .stall_out(Tile_X02_Y0C_stall_out),
    .tile_id(Tile_X02_Y0C_tile_id_in)
);
mantle_wire__typeBit9 Tile_X02_Y0C_hi (
    .in(Tile_X02_Y0C_hi_unq1),
    .out(Tile_X02_Y0C_hi_out)
);
mantle_wire__typeBit8 Tile_X02_Y0C_lo (
    .in(Tile_X02_Y0C_lo_unq1),
    .out(Tile_X02_Y0C_lo_out)
);
wire [15:0] Tile_X02_Y0C_tile_id_out;
assign Tile_X02_Y0C_tile_id_out = {Tile_X02_Y0C_lo_out[7],Tile_X02_Y0C_lo_out[7:6],Tile_X02_Y0C_lo_out[6:5],Tile_X02_Y0C_lo_out[5],Tile_X02_Y0C_hi_out[5],Tile_X02_Y0C_lo_out[4:3],Tile_X02_Y0C_lo_out[3:2],Tile_X02_Y0C_lo_out[2],Tile_X02_Y0C_hi_out[2:1],Tile_X02_Y0C_lo_out[0],Tile_X02_Y0C_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X02_Y0C_tile_id (
    .in(Tile_X02_Y0C_tile_id_in),
    .out(Tile_X02_Y0C_tile_id_out)
);
Tile_PE Tile_X02_Y0D (
    .SB_T0_EAST_SB_IN_B1(Tile_X03_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X03_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X02_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X02_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X02_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X02_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X01_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X01_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X02_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X02_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X03_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X03_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X02_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X02_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X02_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X02_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X01_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X01_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X02_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X02_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X03_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X03_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X02_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X02_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X02_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X02_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X01_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X01_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X02_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X02_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X03_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X03_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X02_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X02_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X02_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X02_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X02_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X02_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X02_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X02_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X01_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X01_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X02_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X02_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X03_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X03_Y0D_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X02_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X02_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X02_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X02_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X02_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X02_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X02_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X02_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X01_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X01_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X02_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X02_Y0D_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y0C_clk_out),
    .clk_out(Tile_X02_Y0D_clk_out),
    .clk_pass_through(Tile_X02_Y0C_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X02_Y0D_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X02_Y0D_clk_pass_through_out_right),
    .config_config_addr(Tile_X02_Y0C_config_out_config_addr),
    .config_config_data(Tile_X02_Y0C_config_out_config_data),
    .config_out_config_addr(Tile_X02_Y0D_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y0D_config_out_config_data),
    .config_out_read(Tile_X02_Y0D_config_out_read),
    .config_out_write(Tile_X02_Y0D_config_out_write),
    .config_read(Tile_X02_Y0C_config_out_read),
    .config_write(Tile_X02_Y0C_config_out_write),
    .hi(Tile_X02_Y0D_hi_unq1),
    .lo(Tile_X02_Y0D_lo_unq1),
    .read_config_data(Tile_X02_Y0D_read_config_data),
    .read_config_data_in(Tile_X02_Y0C_read_config_data),
    .reset(Tile_X02_Y0C_reset_out),
    .reset_out(Tile_X02_Y0D_reset_out),
    .stall(Tile_X02_Y0C_stall_out),
    .stall_out(Tile_X02_Y0D_stall_out),
    .tile_id(Tile_X02_Y0D_tile_id_in)
);
mantle_wire__typeBit9 Tile_X02_Y0D_hi (
    .in(Tile_X02_Y0D_hi_unq1),
    .out(Tile_X02_Y0D_hi_out)
);
mantle_wire__typeBit8 Tile_X02_Y0D_lo (
    .in(Tile_X02_Y0D_lo_unq1),
    .out(Tile_X02_Y0D_lo_out)
);
wire [15:0] Tile_X02_Y0D_tile_id_out;
assign Tile_X02_Y0D_tile_id_out = {Tile_X02_Y0D_lo_out[7],Tile_X02_Y0D_lo_out[7:6],Tile_X02_Y0D_lo_out[6:5],Tile_X02_Y0D_lo_out[5],Tile_X02_Y0D_hi_out[5],Tile_X02_Y0D_lo_out[4:3],Tile_X02_Y0D_lo_out[3:2],Tile_X02_Y0D_lo_out[2],Tile_X02_Y0D_hi_out[2:1],Tile_X02_Y0D_lo_out[0],Tile_X02_Y0D_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X02_Y0D_tile_id (
    .in(Tile_X02_Y0D_tile_id_in),
    .out(Tile_X02_Y0D_tile_id_out)
);
Tile_PE Tile_X02_Y0E (
    .SB_T0_EAST_SB_IN_B1(Tile_X03_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X03_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X02_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X02_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X02_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X02_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X01_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X01_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X02_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X02_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X03_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X03_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X02_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X02_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X02_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X02_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X01_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X01_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X02_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X02_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X03_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X03_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X02_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X02_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X02_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X02_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X01_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X01_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X02_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X02_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X03_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X03_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X02_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X02_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X02_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X02_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X02_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X02_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X02_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X02_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X01_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X01_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X02_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X02_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X03_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X03_Y0E_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X02_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X02_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X02_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X02_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X02_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X02_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X02_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X02_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X01_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X01_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X02_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X02_Y0E_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y0D_clk_out),
    .clk_out(Tile_X02_Y0E_clk_out),
    .clk_pass_through(Tile_X02_Y0D_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X02_Y0E_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X02_Y0E_clk_pass_through_out_right),
    .config_config_addr(Tile_X02_Y0D_config_out_config_addr),
    .config_config_data(Tile_X02_Y0D_config_out_config_data),
    .config_out_config_addr(Tile_X02_Y0E_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y0E_config_out_config_data),
    .config_out_read(Tile_X02_Y0E_config_out_read),
    .config_out_write(Tile_X02_Y0E_config_out_write),
    .config_read(Tile_X02_Y0D_config_out_read),
    .config_write(Tile_X02_Y0D_config_out_write),
    .hi(Tile_X02_Y0E_hi_unq1),
    .lo(Tile_X02_Y0E_lo_unq1),
    .read_config_data(Tile_X02_Y0E_read_config_data),
    .read_config_data_in(Tile_X02_Y0D_read_config_data),
    .reset(Tile_X02_Y0D_reset_out),
    .reset_out(Tile_X02_Y0E_reset_out),
    .stall(Tile_X02_Y0D_stall_out),
    .stall_out(Tile_X02_Y0E_stall_out),
    .tile_id(Tile_X02_Y0E_tile_id_in)
);
mantle_wire__typeBit9 Tile_X02_Y0E_hi (
    .in(Tile_X02_Y0E_hi_unq1),
    .out(Tile_X02_Y0E_hi_out)
);
mantle_wire__typeBit8 Tile_X02_Y0E_lo (
    .in(Tile_X02_Y0E_lo_unq1),
    .out(Tile_X02_Y0E_lo_out)
);
wire [15:0] Tile_X02_Y0E_tile_id_out;
assign Tile_X02_Y0E_tile_id_out = {Tile_X02_Y0E_lo_out[7],Tile_X02_Y0E_lo_out[7:6],Tile_X02_Y0E_lo_out[6:5],Tile_X02_Y0E_lo_out[5],Tile_X02_Y0E_hi_out[5],Tile_X02_Y0E_lo_out[4:3],Tile_X02_Y0E_lo_out[3:2],Tile_X02_Y0E_lo_out[2],Tile_X02_Y0E_hi_out[2:1],Tile_X02_Y0E_hi_out[1],Tile_X02_Y0E_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X02_Y0E_tile_id (
    .in(Tile_X02_Y0E_tile_id_in),
    .out(Tile_X02_Y0E_tile_id_out)
);
Tile_PE Tile_X02_Y0F (
    .SB_T0_EAST_SB_IN_B1(Tile_X03_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X03_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X02_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X02_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X02_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X02_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X02_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X02_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X01_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X01_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X02_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X02_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X03_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X03_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X02_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X02_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X02_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X02_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X02_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X02_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X01_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X01_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X02_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X02_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X03_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X03_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X02_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X02_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X02_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X02_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X02_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X02_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X01_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X01_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X02_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X02_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X03_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X03_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X02_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X02_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X02_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X02_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X02_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X02_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X02_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X02_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X01_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X01_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X02_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X02_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X03_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X03_Y0F_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X02_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X02_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X02_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X02_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X02_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X02_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X02_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X02_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X01_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X01_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X02_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X02_Y0F_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y0E_clk_out),
    .clk_out(Tile_X02_Y0F_clk_out),
    .clk_pass_through(Tile_X02_Y0E_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X02_Y0F_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X02_Y0F_clk_pass_through_out_right),
    .config_config_addr(Tile_X02_Y0E_config_out_config_addr),
    .config_config_data(Tile_X02_Y0E_config_out_config_data),
    .config_out_config_addr(Tile_X02_Y0F_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y0F_config_out_config_data),
    .config_out_read(Tile_X02_Y0F_config_out_read),
    .config_out_write(Tile_X02_Y0F_config_out_write),
    .config_read(Tile_X02_Y0E_config_out_read),
    .config_write(Tile_X02_Y0E_config_out_write),
    .hi(Tile_X02_Y0F_hi_unq1),
    .lo(Tile_X02_Y0F_lo_unq1),
    .read_config_data(Tile_X02_Y0F_read_config_data),
    .read_config_data_in(Tile_X02_Y0E_read_config_data),
    .reset(Tile_X02_Y0E_reset_out),
    .reset_out(Tile_X02_Y0F_reset_out),
    .stall(Tile_X02_Y0E_stall_out),
    .stall_out(Tile_X02_Y0F_stall_out),
    .tile_id(Tile_X02_Y0F_tile_id_in)
);
mantle_wire__typeBit9 Tile_X02_Y0F_hi (
    .in(Tile_X02_Y0F_hi_unq1),
    .out(Tile_X02_Y0F_hi_out)
);
mantle_wire__typeBit8 Tile_X02_Y0F_lo (
    .in(Tile_X02_Y0F_lo_unq1),
    .out(Tile_X02_Y0F_lo_out)
);
wire [15:0] Tile_X02_Y0F_tile_id_out;
assign Tile_X02_Y0F_tile_id_out = {Tile_X02_Y0F_lo_out[7],Tile_X02_Y0F_lo_out[7:6],Tile_X02_Y0F_lo_out[6:5],Tile_X02_Y0F_lo_out[5],Tile_X02_Y0F_hi_out[5],Tile_X02_Y0F_lo_out[4:3],Tile_X02_Y0F_lo_out[3:2],Tile_X02_Y0F_lo_out[2],Tile_X02_Y0F_hi_out[2:1],Tile_X02_Y0F_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X02_Y0F_tile_id (
    .in(Tile_X02_Y0F_tile_id_in),
    .out(Tile_X02_Y0F_tile_id_out)
);
Tile_PE Tile_X02_Y10 (
    .SB_T0_EAST_SB_IN_B1(Tile_X03_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X03_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X02_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X02_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X02_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X02_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X02_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X02_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T0_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X02_Y10_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X02_Y10_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X01_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X01_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X02_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X02_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X03_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X03_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X02_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X02_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X02_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X02_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X02_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X02_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T1_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X02_Y10_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X02_Y10_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X01_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X01_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X02_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X02_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X03_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X03_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X02_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X02_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X02_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X02_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X02_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X02_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T2_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X02_Y10_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X02_Y10_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X01_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X01_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X02_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X02_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X03_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X03_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X02_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X02_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X02_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X02_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X02_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X02_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T3_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X02_Y10_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X02_Y10_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X01_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X01_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X02_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X02_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X03_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X03_Y10_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X02_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X02_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X02_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X02_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X02_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X02_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T4_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X02_Y10_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X02_Y10_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X01_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X01_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X02_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X02_Y10_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y0F_clk_out),
    .clk_out(Tile_X02_Y10_clk_out),
    .clk_pass_through(Tile_X02_Y0F_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X02_Y10_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X02_Y10_clk_pass_through_out_right),
    .config_config_addr(Tile_X02_Y0F_config_out_config_addr),
    .config_config_data(Tile_X02_Y0F_config_out_config_data),
    .config_out_config_addr(Tile_X02_Y10_config_out_config_addr),
    .config_out_config_data(Tile_X02_Y10_config_out_config_data),
    .config_out_read(Tile_X02_Y10_config_out_read),
    .config_out_write(Tile_X02_Y10_config_out_write),
    .config_read(Tile_X02_Y0F_config_out_read),
    .config_write(Tile_X02_Y0F_config_out_write),
    .hi(Tile_X02_Y10_hi),
    .lo(Tile_X02_Y10_lo_unq1),
    .read_config_data(Tile_X02_Y10_read_config_data),
    .read_config_data_in(Tile_X02_Y0F_read_config_data),
    .reset(Tile_X02_Y0F_reset_out),
    .reset_out(Tile_X02_Y10_reset_out),
    .stall(Tile_X02_Y0F_stall_out),
    .stall_out(Tile_X02_Y10_stall_out),
    .tile_id(Tile_X02_Y10_tile_id_in)
);
mantle_wire__typeBit8 Tile_X02_Y10_lo (
    .in(Tile_X02_Y10_lo_unq1),
    .out(Tile_X02_Y10_lo_out)
);
wire [15:0] Tile_X02_Y10_tile_id_out;
assign Tile_X02_Y10_tile_id_out = {Tile_X02_Y10_lo_out[7],Tile_X02_Y10_lo_out[7:6],Tile_X02_Y10_lo_out[6:5],Tile_X02_Y10_lo_out[5],Tile_X02_Y10_hi[5],Tile_X02_Y10_lo_out[4:3],Tile_X02_Y10_lo_out[3:2],Tile_X02_Y10_hi[2],Tile_X02_Y10_lo_out[1],Tile_X02_Y10_lo_out[1:0],Tile_X02_Y10_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X02_Y10_tile_id (
    .in(Tile_X02_Y10_tile_id_in),
    .out(Tile_X02_Y10_tile_id_out)
);
wire [15:0] Tile_X03_Y00_tile_id;
assign Tile_X03_Y00_tile_id = {Tile_X03_Y00_lo[7],Tile_X03_Y00_lo[7:6],Tile_X03_Y00_lo[6:5],Tile_X03_Y00_lo[5],Tile_X03_Y00_hi[5:4],Tile_X03_Y00_lo[3],Tile_X03_Y00_lo[3:2],Tile_X03_Y00_lo[2:1],Tile_X03_Y00_lo[1:0],Tile_X03_Y00_lo[0]};
Tile_io_core Tile_X03_Y00 (
    .tile_id(Tile_X03_Y00_tile_id),
    .glb2io_1(glb2io_1_X03_Y00),
    .f2io_1(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B1),
    .io2glb_1(Tile_X03_Y00_io2glb_1),
    .io2f_1(Tile_X03_Y00_io2f_1),
    .glb2io_16(glb2io_16_X03_Y00),
    .f2io_16(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B16),
    .io2glb_16(Tile_X03_Y00_io2glb_16),
    .io2f_16(Tile_X03_Y00_io2f_16),
    .hi(Tile_X03_Y00_hi),
    .lo(Tile_X03_Y00_lo)
);
Tile_MemCore Tile_X03_Y01 (
    .SB_T0_EAST_SB_IN_B1(Tile_X04_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X04_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X03_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X03_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X03_Y00_io2f_1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X03_Y00_io2f_16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y01_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X02_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X03_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X04_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X04_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X03_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X03_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X03_Y00_io2f_1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X03_Y00_io2f_16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y01_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X02_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X03_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X04_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X04_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X03_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X03_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X03_Y00_io2f_1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X03_Y00_io2f_16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y01_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X02_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X03_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X04_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X04_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X03_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X03_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X03_Y00_io2f_1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X03_Y00_io2f_16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y01_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X03_Y01_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X02_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X02_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X03_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X03_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X04_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X04_Y01_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X03_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X03_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X03_Y00_io2f_1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X03_Y00_io2f_16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y01_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X03_Y01_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X02_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X02_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X03_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X03_Y01_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y01_clk_pass_through_out_right),
    .clk_out(Tile_X03_Y01_clk_out),
    .config_config_addr(config_3_config_addr),
    .config_config_data(config_3_config_data),
    .config_out_config_addr(Tile_X03_Y01_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y01_config_out_config_data),
    .config_out_read(Tile_X03_Y01_config_out_read),
    .config_out_write(Tile_X03_Y01_config_out_write),
    .config_read(config_3_read),
    .config_write(config_3_write),
    .hi(Tile_X03_Y01_hi_unq1),
    .lo(Tile_X03_Y01_lo_unq1),
    .read_config_data(Tile_X03_Y01_read_config_data),
    .read_config_data_in(const_0_32_out),
    .reset(reset),
    .reset_out(Tile_X03_Y01_reset_out),
    .stall(stall[3]),
    .stall_out(Tile_X03_Y01_stall_out),
    .tile_id(Tile_X03_Y01_tile_id_in)
);
mantle_wire__typeBit9 Tile_X03_Y01_hi (
    .in(Tile_X03_Y01_hi_unq1),
    .out(Tile_X03_Y01_hi_out)
);
mantle_wire__typeBit8 Tile_X03_Y01_lo (
    .in(Tile_X03_Y01_lo_unq1),
    .out(Tile_X03_Y01_lo_out)
);
wire [15:0] Tile_X03_Y01_tile_id_out;
assign Tile_X03_Y01_tile_id_out = {Tile_X03_Y01_lo_out[7],Tile_X03_Y01_lo_out[7:6],Tile_X03_Y01_lo_out[6:5],Tile_X03_Y01_lo_out[5],Tile_X03_Y01_hi_out[5:4],Tile_X03_Y01_lo_out[3],Tile_X03_Y01_lo_out[3:2],Tile_X03_Y01_lo_out[2:1],Tile_X03_Y01_lo_out[1:0],Tile_X03_Y01_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X03_Y01_tile_id (
    .in(Tile_X03_Y01_tile_id_in),
    .out(Tile_X03_Y01_tile_id_out)
);
Tile_MemCore Tile_X03_Y02 (
    .SB_T0_EAST_SB_IN_B1(Tile_X04_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X04_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X03_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X03_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X03_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X02_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X03_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X04_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X04_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X03_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X03_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X03_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X02_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X03_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X04_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X04_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X03_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X03_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X03_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X02_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X03_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X04_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X04_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X03_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X03_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X03_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X03_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X02_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X02_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X03_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X03_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X04_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X04_Y02_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X03_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X03_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X03_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X03_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X02_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X02_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X03_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X03_Y02_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y02_clk_pass_through_out_right),
    .clk_out(Tile_X03_Y02_clk_out),
    .config_config_addr(Tile_X03_Y01_config_out_config_addr),
    .config_config_data(Tile_X03_Y01_config_out_config_data),
    .config_out_config_addr(Tile_X03_Y02_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y02_config_out_config_data),
    .config_out_read(Tile_X03_Y02_config_out_read),
    .config_out_write(Tile_X03_Y02_config_out_write),
    .config_read(Tile_X03_Y01_config_out_read),
    .config_write(Tile_X03_Y01_config_out_write),
    .hi(Tile_X03_Y02_hi_unq1),
    .lo(Tile_X03_Y02_lo_unq1),
    .read_config_data(Tile_X03_Y02_read_config_data),
    .read_config_data_in(Tile_X03_Y01_read_config_data),
    .reset(Tile_X03_Y01_reset_out),
    .reset_out(Tile_X03_Y02_reset_out),
    .stall(Tile_X03_Y01_stall_out),
    .stall_out(Tile_X03_Y02_stall_out),
    .tile_id(Tile_X03_Y02_tile_id_in)
);
mantle_wire__typeBit9 Tile_X03_Y02_hi (
    .in(Tile_X03_Y02_hi_unq1),
    .out(Tile_X03_Y02_hi_out)
);
mantle_wire__typeBit8 Tile_X03_Y02_lo (
    .in(Tile_X03_Y02_lo_unq1),
    .out(Tile_X03_Y02_lo_out)
);
wire [15:0] Tile_X03_Y02_tile_id_out;
assign Tile_X03_Y02_tile_id_out = {Tile_X03_Y02_lo_out[7],Tile_X03_Y02_lo_out[7:6],Tile_X03_Y02_lo_out[6:5],Tile_X03_Y02_lo_out[5],Tile_X03_Y02_hi_out[5:4],Tile_X03_Y02_lo_out[3],Tile_X03_Y02_lo_out[3:2],Tile_X03_Y02_lo_out[2:1],Tile_X03_Y02_lo_out[1],Tile_X03_Y02_hi_out[1],Tile_X03_Y02_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X03_Y02_tile_id (
    .in(Tile_X03_Y02_tile_id_in),
    .out(Tile_X03_Y02_tile_id_out)
);
Tile_MemCore Tile_X03_Y03 (
    .SB_T0_EAST_SB_IN_B1(Tile_X04_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X04_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X03_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X03_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X03_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X02_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X03_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X04_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X04_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X03_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X03_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X03_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X02_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X03_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X04_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X04_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X03_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X03_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X03_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X02_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X03_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X04_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X04_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X03_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X03_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X03_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X03_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X02_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X02_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X03_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X03_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X04_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X04_Y03_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X03_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X03_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X03_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X03_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X02_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X02_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X03_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X03_Y03_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y03_clk_pass_through_out_right),
    .clk_out(Tile_X03_Y03_clk_out),
    .config_config_addr(Tile_X03_Y02_config_out_config_addr),
    .config_config_data(Tile_X03_Y02_config_out_config_data),
    .config_out_config_addr(Tile_X03_Y03_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y03_config_out_config_data),
    .config_out_read(Tile_X03_Y03_config_out_read),
    .config_out_write(Tile_X03_Y03_config_out_write),
    .config_read(Tile_X03_Y02_config_out_read),
    .config_write(Tile_X03_Y02_config_out_write),
    .hi(Tile_X03_Y03_hi_unq1),
    .lo(Tile_X03_Y03_lo_unq1),
    .read_config_data(Tile_X03_Y03_read_config_data),
    .read_config_data_in(Tile_X03_Y02_read_config_data),
    .reset(Tile_X03_Y02_reset_out),
    .reset_out(Tile_X03_Y03_reset_out),
    .stall(Tile_X03_Y02_stall_out),
    .stall_out(Tile_X03_Y03_stall_out),
    .tile_id(Tile_X03_Y03_tile_id_in)
);
mantle_wire__typeBit9 Tile_X03_Y03_hi (
    .in(Tile_X03_Y03_hi_unq1),
    .out(Tile_X03_Y03_hi_out)
);
mantle_wire__typeBit8 Tile_X03_Y03_lo (
    .in(Tile_X03_Y03_lo_unq1),
    .out(Tile_X03_Y03_lo_out)
);
wire [15:0] Tile_X03_Y03_tile_id_out;
assign Tile_X03_Y03_tile_id_out = {Tile_X03_Y03_lo_out[7],Tile_X03_Y03_lo_out[7:6],Tile_X03_Y03_lo_out[6:5],Tile_X03_Y03_lo_out[5],Tile_X03_Y03_hi_out[5:4],Tile_X03_Y03_lo_out[3],Tile_X03_Y03_lo_out[3:2],Tile_X03_Y03_lo_out[2:1],Tile_X03_Y03_lo_out[1],Tile_X03_Y03_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X03_Y03_tile_id (
    .in(Tile_X03_Y03_tile_id_in),
    .out(Tile_X03_Y03_tile_id_out)
);
Tile_MemCore Tile_X03_Y04 (
    .SB_T0_EAST_SB_IN_B1(Tile_X04_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X04_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X03_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X03_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X03_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X02_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X03_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X04_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X04_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X03_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X03_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X03_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X02_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X03_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X04_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X04_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X03_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X03_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X03_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X02_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X03_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X04_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X04_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X03_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X03_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X03_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X03_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X03_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X03_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X02_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X02_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X03_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X03_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X04_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X04_Y04_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X03_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X03_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X03_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X03_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X03_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X03_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X02_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X02_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X03_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X03_Y04_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y04_clk_pass_through_out_right),
    .clk_out(Tile_X03_Y04_clk_out),
    .config_config_addr(Tile_X03_Y03_config_out_config_addr),
    .config_config_data(Tile_X03_Y03_config_out_config_data),
    .config_out_config_addr(Tile_X03_Y04_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y04_config_out_config_data),
    .config_out_read(Tile_X03_Y04_config_out_read),
    .config_out_write(Tile_X03_Y04_config_out_write),
    .config_read(Tile_X03_Y03_config_out_read),
    .config_write(Tile_X03_Y03_config_out_write),
    .hi(Tile_X03_Y04_hi_unq1),
    .lo(Tile_X03_Y04_lo_unq1),
    .read_config_data(Tile_X03_Y04_read_config_data),
    .read_config_data_in(Tile_X03_Y03_read_config_data),
    .reset(Tile_X03_Y03_reset_out),
    .reset_out(Tile_X03_Y04_reset_out),
    .stall(Tile_X03_Y03_stall_out),
    .stall_out(Tile_X03_Y04_stall_out),
    .tile_id(Tile_X03_Y04_tile_id_in)
);
mantle_wire__typeBit9 Tile_X03_Y04_hi (
    .in(Tile_X03_Y04_hi_unq1),
    .out(Tile_X03_Y04_hi_out)
);
mantle_wire__typeBit8 Tile_X03_Y04_lo (
    .in(Tile_X03_Y04_lo_unq1),
    .out(Tile_X03_Y04_lo_out)
);
wire [15:0] Tile_X03_Y04_tile_id_out;
assign Tile_X03_Y04_tile_id_out = {Tile_X03_Y04_lo_out[7],Tile_X03_Y04_lo_out[7:6],Tile_X03_Y04_lo_out[6:5],Tile_X03_Y04_lo_out[5],Tile_X03_Y04_hi_out[5:4],Tile_X03_Y04_lo_out[3],Tile_X03_Y04_lo_out[3:2],Tile_X03_Y04_lo_out[2:1],Tile_X03_Y04_hi_out[1],Tile_X03_Y04_lo_out[0],Tile_X03_Y04_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X03_Y04_tile_id (
    .in(Tile_X03_Y04_tile_id_in),
    .out(Tile_X03_Y04_tile_id_out)
);
Tile_MemCore Tile_X03_Y05 (
    .SB_T0_EAST_SB_IN_B1(Tile_X04_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X04_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X03_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X03_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X03_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X02_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X02_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X03_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X03_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X04_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X04_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X03_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X03_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X03_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X02_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X02_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X03_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X03_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X04_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X04_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X03_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X03_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X03_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X02_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X02_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X03_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X03_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X04_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X04_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X03_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X03_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X03_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X03_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X03_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X03_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X03_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X02_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X02_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X03_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X03_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X04_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X04_Y05_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X03_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X03_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X03_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X03_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X03_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X03_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X03_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X02_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X02_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X03_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X03_Y05_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y05_clk_pass_through_out_right),
    .clk_out(Tile_X03_Y05_clk_out),
    .config_config_addr(Tile_X03_Y04_config_out_config_addr),
    .config_config_data(Tile_X03_Y04_config_out_config_data),
    .config_out_config_addr(Tile_X03_Y05_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y05_config_out_config_data),
    .config_out_read(Tile_X03_Y05_config_out_read),
    .config_out_write(Tile_X03_Y05_config_out_write),
    .config_read(Tile_X03_Y04_config_out_read),
    .config_write(Tile_X03_Y04_config_out_write),
    .hi(Tile_X03_Y05_hi_unq1),
    .lo(Tile_X03_Y05_lo_unq1),
    .read_config_data(Tile_X03_Y05_read_config_data),
    .read_config_data_in(Tile_X03_Y04_read_config_data),
    .reset(Tile_X03_Y04_reset_out),
    .reset_out(Tile_X03_Y05_reset_out),
    .stall(Tile_X03_Y04_stall_out),
    .stall_out(Tile_X03_Y05_stall_out),
    .tile_id(Tile_X03_Y05_tile_id_in)
);
mantle_wire__typeBit9 Tile_X03_Y05_hi (
    .in(Tile_X03_Y05_hi_unq1),
    .out(Tile_X03_Y05_hi_out)
);
mantle_wire__typeBit8 Tile_X03_Y05_lo (
    .in(Tile_X03_Y05_lo_unq1),
    .out(Tile_X03_Y05_lo_out)
);
wire [15:0] Tile_X03_Y05_tile_id_out;
assign Tile_X03_Y05_tile_id_out = {Tile_X03_Y05_lo_out[7],Tile_X03_Y05_lo_out[7:6],Tile_X03_Y05_lo_out[6:5],Tile_X03_Y05_lo_out[5],Tile_X03_Y05_hi_out[5:4],Tile_X03_Y05_lo_out[3],Tile_X03_Y05_lo_out[3:2],Tile_X03_Y05_lo_out[2:1],Tile_X03_Y05_hi_out[1],Tile_X03_Y05_lo_out[0],Tile_X03_Y05_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X03_Y05_tile_id (
    .in(Tile_X03_Y05_tile_id_in),
    .out(Tile_X03_Y05_tile_id_out)
);
Tile_MemCore Tile_X03_Y06 (
    .SB_T0_EAST_SB_IN_B1(Tile_X04_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X04_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X03_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X03_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X03_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X03_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X02_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X02_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X03_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X03_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X04_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X04_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X03_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X03_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X03_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X03_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X02_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X02_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X03_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X03_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X04_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X04_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X03_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X03_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X03_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X03_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X02_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X02_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X03_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X03_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X04_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X04_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X03_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X03_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X03_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X03_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X03_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X03_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X03_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X03_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X02_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X02_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X03_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X03_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X04_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X04_Y06_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X03_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X03_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X03_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X03_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X03_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X03_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X03_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X03_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X02_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X02_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X03_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X03_Y06_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y06_clk_pass_through_out_right),
    .clk_out(Tile_X03_Y06_clk_out),
    .config_config_addr(Tile_X03_Y05_config_out_config_addr),
    .config_config_data(Tile_X03_Y05_config_out_config_data),
    .config_out_config_addr(Tile_X03_Y06_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y06_config_out_config_data),
    .config_out_read(Tile_X03_Y06_config_out_read),
    .config_out_write(Tile_X03_Y06_config_out_write),
    .config_read(Tile_X03_Y05_config_out_read),
    .config_write(Tile_X03_Y05_config_out_write),
    .hi(Tile_X03_Y06_hi_unq1),
    .lo(Tile_X03_Y06_lo_unq1),
    .read_config_data(Tile_X03_Y06_read_config_data),
    .read_config_data_in(Tile_X03_Y05_read_config_data),
    .reset(Tile_X03_Y05_reset_out),
    .reset_out(Tile_X03_Y06_reset_out),
    .stall(Tile_X03_Y05_stall_out),
    .stall_out(Tile_X03_Y06_stall_out),
    .tile_id(Tile_X03_Y06_tile_id_in)
);
mantle_wire__typeBit9 Tile_X03_Y06_hi (
    .in(Tile_X03_Y06_hi_unq1),
    .out(Tile_X03_Y06_hi_out)
);
mantle_wire__typeBit8 Tile_X03_Y06_lo (
    .in(Tile_X03_Y06_lo_unq1),
    .out(Tile_X03_Y06_lo_out)
);
wire [15:0] Tile_X03_Y06_tile_id_out;
assign Tile_X03_Y06_tile_id_out = {Tile_X03_Y06_lo_out[7],Tile_X03_Y06_lo_out[7:6],Tile_X03_Y06_lo_out[6:5],Tile_X03_Y06_lo_out[5],Tile_X03_Y06_hi_out[5:4],Tile_X03_Y06_lo_out[3],Tile_X03_Y06_lo_out[3:2],Tile_X03_Y06_lo_out[2:1],Tile_X03_Y06_hi_out[1],Tile_X03_Y06_hi_out[1],Tile_X03_Y06_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X03_Y06_tile_id (
    .in(Tile_X03_Y06_tile_id_in),
    .out(Tile_X03_Y06_tile_id_out)
);
Tile_MemCore Tile_X03_Y07 (
    .SB_T0_EAST_SB_IN_B1(Tile_X04_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X04_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X03_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X03_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X03_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X03_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X02_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X02_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X03_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X03_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X04_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X04_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X03_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X03_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X03_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X03_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X02_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X02_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X03_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X03_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X04_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X04_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X03_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X03_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X03_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X03_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X02_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X02_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X03_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X03_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X04_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X04_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X03_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X03_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X03_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X03_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X03_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X03_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X03_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X03_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X02_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X02_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X03_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X03_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X04_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X04_Y07_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X03_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X03_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X03_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X03_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X03_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X03_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X03_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X03_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X02_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X02_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X03_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X03_Y07_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y07_clk_pass_through_out_right),
    .clk_out(Tile_X03_Y07_clk_out),
    .config_config_addr(Tile_X03_Y06_config_out_config_addr),
    .config_config_data(Tile_X03_Y06_config_out_config_data),
    .config_out_config_addr(Tile_X03_Y07_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y07_config_out_config_data),
    .config_out_read(Tile_X03_Y07_config_out_read),
    .config_out_write(Tile_X03_Y07_config_out_write),
    .config_read(Tile_X03_Y06_config_out_read),
    .config_write(Tile_X03_Y06_config_out_write),
    .hi(Tile_X03_Y07_hi_unq1),
    .lo(Tile_X03_Y07_lo_unq1),
    .read_config_data(Tile_X03_Y07_read_config_data),
    .read_config_data_in(Tile_X03_Y06_read_config_data),
    .reset(Tile_X03_Y06_reset_out),
    .reset_out(Tile_X03_Y07_reset_out),
    .stall(Tile_X03_Y06_stall_out),
    .stall_out(Tile_X03_Y07_stall_out),
    .tile_id(Tile_X03_Y07_tile_id_in)
);
mantle_wire__typeBit9 Tile_X03_Y07_hi (
    .in(Tile_X03_Y07_hi_unq1),
    .out(Tile_X03_Y07_hi_out)
);
mantle_wire__typeBit8 Tile_X03_Y07_lo (
    .in(Tile_X03_Y07_lo_unq1),
    .out(Tile_X03_Y07_lo_out)
);
wire [15:0] Tile_X03_Y07_tile_id_out;
assign Tile_X03_Y07_tile_id_out = {Tile_X03_Y07_lo_out[7],Tile_X03_Y07_lo_out[7:6],Tile_X03_Y07_lo_out[6:5],Tile_X03_Y07_lo_out[5],Tile_X03_Y07_hi_out[5:4],Tile_X03_Y07_lo_out[3],Tile_X03_Y07_lo_out[3:2],Tile_X03_Y07_lo_out[2:1],Tile_X03_Y07_hi_out[1],Tile_X03_Y07_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X03_Y07_tile_id (
    .in(Tile_X03_Y07_tile_id_in),
    .out(Tile_X03_Y07_tile_id_out)
);
Tile_MemCore Tile_X03_Y08 (
    .SB_T0_EAST_SB_IN_B1(Tile_X04_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X04_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X03_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X03_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X03_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X03_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X02_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X02_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X03_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X03_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X04_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X04_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X03_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X03_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X03_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X03_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X02_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X02_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X03_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X03_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X04_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X04_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X03_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X03_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X03_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X03_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X02_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X02_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X03_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X03_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X04_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X04_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X03_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X03_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X03_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X03_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X03_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X03_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X03_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X03_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X02_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X02_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X03_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X03_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X04_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X04_Y08_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X03_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X03_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X03_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X03_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X03_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X03_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X03_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X03_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X02_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X02_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X03_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X03_Y08_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y08_clk_pass_through_out_right),
    .clk_out(Tile_X03_Y08_clk_out),
    .config_config_addr(Tile_X03_Y07_config_out_config_addr),
    .config_config_data(Tile_X03_Y07_config_out_config_data),
    .config_out_config_addr(Tile_X03_Y08_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y08_config_out_config_data),
    .config_out_read(Tile_X03_Y08_config_out_read),
    .config_out_write(Tile_X03_Y08_config_out_write),
    .config_read(Tile_X03_Y07_config_out_read),
    .config_write(Tile_X03_Y07_config_out_write),
    .hi(Tile_X03_Y08_hi_unq1),
    .lo(Tile_X03_Y08_lo_unq1),
    .read_config_data(Tile_X03_Y08_read_config_data),
    .read_config_data_in(Tile_X03_Y07_read_config_data),
    .reset(Tile_X03_Y07_reset_out),
    .reset_out(Tile_X03_Y08_reset_out),
    .stall(Tile_X03_Y07_stall_out),
    .stall_out(Tile_X03_Y08_stall_out),
    .tile_id(Tile_X03_Y08_tile_id_in)
);
mantle_wire__typeBit9 Tile_X03_Y08_hi (
    .in(Tile_X03_Y08_hi_unq1),
    .out(Tile_X03_Y08_hi_out)
);
mantle_wire__typeBit8 Tile_X03_Y08_lo (
    .in(Tile_X03_Y08_lo_unq1),
    .out(Tile_X03_Y08_lo_out)
);
wire [15:0] Tile_X03_Y08_tile_id_out;
assign Tile_X03_Y08_tile_id_out = {Tile_X03_Y08_lo_out[7],Tile_X03_Y08_lo_out[7:6],Tile_X03_Y08_lo_out[6:5],Tile_X03_Y08_lo_out[5],Tile_X03_Y08_hi_out[5:4],Tile_X03_Y08_lo_out[3],Tile_X03_Y08_lo_out[3:2],Tile_X03_Y08_lo_out[2],Tile_X03_Y08_hi_out[2],Tile_X03_Y08_lo_out[1:0],Tile_X03_Y08_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X03_Y08_tile_id (
    .in(Tile_X03_Y08_tile_id_in),
    .out(Tile_X03_Y08_tile_id_out)
);
Tile_MemCore Tile_X03_Y09 (
    .SB_T0_EAST_SB_IN_B1(Tile_X04_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X04_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X03_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X03_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X03_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X03_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X02_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X02_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X03_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X03_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X04_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X04_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X03_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X03_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X03_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X03_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X02_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X02_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X03_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X03_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X04_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X04_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X03_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X03_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X03_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X03_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X02_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X02_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X03_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X03_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X04_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X04_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X03_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X03_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X03_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X03_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X03_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X03_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X03_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X03_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X02_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X02_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X03_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X03_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X04_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X04_Y09_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X03_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X03_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X03_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X03_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X03_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X03_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X03_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X03_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X02_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X02_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X03_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X03_Y09_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y09_clk_pass_through_out_right),
    .clk_out(Tile_X03_Y09_clk_out),
    .config_config_addr(ConfigPipeStage_inst3_config_out_config_addr),
    .config_config_data(ConfigPipeStage_inst3_config_out_config_data),
    .config_out_config_addr(Tile_X03_Y09_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y09_config_out_config_data),
    .config_out_read(Tile_X03_Y09_config_out_read),
    .config_out_write(Tile_X03_Y09_config_out_write),
    .config_read(ConfigPipeStage_inst3_config_out_read),
    .config_write(ConfigPipeStage_inst3_config_out_write),
    .hi(Tile_X03_Y09_hi_unq1),
    .lo(Tile_X03_Y09_lo_unq1),
    .read_config_data(Tile_X03_Y09_read_config_data),
    .read_config_data_in(Tile_X03_Y08_read_config_data),
    .reset(Tile_X03_Y08_reset_out),
    .reset_out(Tile_X03_Y09_reset_out),
    .stall(Tile_X03_Y08_stall_out),
    .stall_out(Tile_X03_Y09_stall_out),
    .tile_id(Tile_X03_Y09_tile_id_in)
);
mantle_wire__typeBit9 Tile_X03_Y09_hi (
    .in(Tile_X03_Y09_hi_unq1),
    .out(Tile_X03_Y09_hi_out)
);
mantle_wire__typeBit8 Tile_X03_Y09_lo (
    .in(Tile_X03_Y09_lo_unq1),
    .out(Tile_X03_Y09_lo_out)
);
wire [15:0] Tile_X03_Y09_tile_id_out;
assign Tile_X03_Y09_tile_id_out = {Tile_X03_Y09_lo_out[7],Tile_X03_Y09_lo_out[7:6],Tile_X03_Y09_lo_out[6:5],Tile_X03_Y09_lo_out[5],Tile_X03_Y09_hi_out[5:4],Tile_X03_Y09_lo_out[3],Tile_X03_Y09_lo_out[3:2],Tile_X03_Y09_lo_out[2],Tile_X03_Y09_hi_out[2],Tile_X03_Y09_lo_out[1:0],Tile_X03_Y09_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X03_Y09_tile_id (
    .in(Tile_X03_Y09_tile_id_in),
    .out(Tile_X03_Y09_tile_id_out)
);
Tile_MemCore Tile_X03_Y0A (
    .SB_T0_EAST_SB_IN_B1(Tile_X04_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X04_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X03_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X03_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X03_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X03_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X02_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X02_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X03_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X03_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X04_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X04_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X03_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X03_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X03_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X03_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X02_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X02_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X03_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X03_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X04_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X04_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X03_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X03_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X03_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X03_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X02_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X02_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X03_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X03_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X04_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X04_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X03_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X03_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X03_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X03_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X03_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X03_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X03_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X03_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X02_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X02_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X03_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X03_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X04_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X04_Y0A_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X03_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X03_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X03_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X03_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X03_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X03_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X03_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X03_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X02_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X02_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X03_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X03_Y0A_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y0A_clk_pass_through_out_right),
    .clk_out(Tile_X03_Y0A_clk_out),
    .config_config_addr(Tile_X03_Y09_config_out_config_addr),
    .config_config_data(Tile_X03_Y09_config_out_config_data),
    .config_out_config_addr(Tile_X03_Y0A_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y0A_config_out_config_data),
    .config_out_read(Tile_X03_Y0A_config_out_read),
    .config_out_write(Tile_X03_Y0A_config_out_write),
    .config_read(Tile_X03_Y09_config_out_read),
    .config_write(Tile_X03_Y09_config_out_write),
    .hi(Tile_X03_Y0A_hi_unq1),
    .lo(Tile_X03_Y0A_lo_unq1),
    .read_config_data(Tile_X03_Y0A_read_config_data),
    .read_config_data_in(Tile_X03_Y09_read_config_data),
    .reset(Tile_X03_Y09_reset_out),
    .reset_out(Tile_X03_Y0A_reset_out),
    .stall(Tile_X03_Y09_stall_out),
    .stall_out(Tile_X03_Y0A_stall_out),
    .tile_id(Tile_X03_Y0A_tile_id_in)
);
mantle_wire__typeBit9 Tile_X03_Y0A_hi (
    .in(Tile_X03_Y0A_hi_unq1),
    .out(Tile_X03_Y0A_hi_out)
);
mantle_wire__typeBit8 Tile_X03_Y0A_lo (
    .in(Tile_X03_Y0A_lo_unq1),
    .out(Tile_X03_Y0A_lo_out)
);
wire [15:0] Tile_X03_Y0A_tile_id_out;
assign Tile_X03_Y0A_tile_id_out = {Tile_X03_Y0A_lo_out[7],Tile_X03_Y0A_lo_out[7:6],Tile_X03_Y0A_lo_out[6:5],Tile_X03_Y0A_lo_out[5],Tile_X03_Y0A_hi_out[5:4],Tile_X03_Y0A_lo_out[3],Tile_X03_Y0A_lo_out[3:2],Tile_X03_Y0A_lo_out[2],Tile_X03_Y0A_hi_out[2],Tile_X03_Y0A_lo_out[1],Tile_X03_Y0A_hi_out[1],Tile_X03_Y0A_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X03_Y0A_tile_id (
    .in(Tile_X03_Y0A_tile_id_in),
    .out(Tile_X03_Y0A_tile_id_out)
);
Tile_MemCore Tile_X03_Y0B (
    .SB_T0_EAST_SB_IN_B1(Tile_X04_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X04_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X03_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X03_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X03_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X03_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X02_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X02_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X03_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X03_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X04_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X04_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X03_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X03_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X03_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X03_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X02_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X02_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X03_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X03_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X04_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X04_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X03_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X03_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X03_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X03_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X02_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X02_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X03_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X03_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X04_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X04_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X03_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X03_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X03_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X03_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X03_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X03_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X03_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X03_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X02_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X02_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X03_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X03_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X04_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X04_Y0B_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X03_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X03_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X03_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X03_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X03_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X03_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X03_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X03_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X02_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X02_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X03_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X03_Y0B_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y0B_clk_pass_through_out_right),
    .clk_out(Tile_X03_Y0B_clk_out),
    .config_config_addr(Tile_X03_Y0A_config_out_config_addr),
    .config_config_data(Tile_X03_Y0A_config_out_config_data),
    .config_out_config_addr(Tile_X03_Y0B_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y0B_config_out_config_data),
    .config_out_read(Tile_X03_Y0B_config_out_read),
    .config_out_write(Tile_X03_Y0B_config_out_write),
    .config_read(Tile_X03_Y0A_config_out_read),
    .config_write(Tile_X03_Y0A_config_out_write),
    .hi(Tile_X03_Y0B_hi_unq1),
    .lo(Tile_X03_Y0B_lo_unq1),
    .read_config_data(Tile_X03_Y0B_read_config_data),
    .read_config_data_in(Tile_X03_Y0A_read_config_data),
    .reset(Tile_X03_Y0A_reset_out),
    .reset_out(Tile_X03_Y0B_reset_out),
    .stall(Tile_X03_Y0A_stall_out),
    .stall_out(Tile_X03_Y0B_stall_out),
    .tile_id(Tile_X03_Y0B_tile_id_in)
);
mantle_wire__typeBit9 Tile_X03_Y0B_hi (
    .in(Tile_X03_Y0B_hi_unq1),
    .out(Tile_X03_Y0B_hi_out)
);
mantle_wire__typeBit8 Tile_X03_Y0B_lo (
    .in(Tile_X03_Y0B_lo_unq1),
    .out(Tile_X03_Y0B_lo_out)
);
wire [15:0] Tile_X03_Y0B_tile_id_out;
assign Tile_X03_Y0B_tile_id_out = {Tile_X03_Y0B_lo_out[7],Tile_X03_Y0B_lo_out[7:6],Tile_X03_Y0B_lo_out[6:5],Tile_X03_Y0B_lo_out[5],Tile_X03_Y0B_hi_out[5:4],Tile_X03_Y0B_lo_out[3],Tile_X03_Y0B_lo_out[3:2],Tile_X03_Y0B_lo_out[2],Tile_X03_Y0B_hi_out[2],Tile_X03_Y0B_lo_out[1],Tile_X03_Y0B_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X03_Y0B_tile_id (
    .in(Tile_X03_Y0B_tile_id_in),
    .out(Tile_X03_Y0B_tile_id_out)
);
Tile_MemCore Tile_X03_Y0C (
    .SB_T0_EAST_SB_IN_B1(Tile_X04_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X04_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X03_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X03_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X03_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X03_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X02_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X02_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X03_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X03_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X04_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X04_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X03_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X03_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X03_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X03_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X02_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X02_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X03_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X03_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X04_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X04_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X03_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X03_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X03_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X03_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X02_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X02_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X03_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X03_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X04_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X04_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X03_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X03_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X03_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X03_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X03_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X03_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X03_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X03_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X02_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X02_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X03_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X03_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X04_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X04_Y0C_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X03_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X03_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X03_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X03_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X03_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X03_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X03_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X03_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X02_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X02_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X03_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X03_Y0C_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y0C_clk_pass_through_out_right),
    .clk_out(Tile_X03_Y0C_clk_out),
    .config_config_addr(Tile_X03_Y0B_config_out_config_addr),
    .config_config_data(Tile_X03_Y0B_config_out_config_data),
    .config_out_config_addr(Tile_X03_Y0C_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y0C_config_out_config_data),
    .config_out_read(Tile_X03_Y0C_config_out_read),
    .config_out_write(Tile_X03_Y0C_config_out_write),
    .config_read(Tile_X03_Y0B_config_out_read),
    .config_write(Tile_X03_Y0B_config_out_write),
    .hi(Tile_X03_Y0C_hi_unq1),
    .lo(Tile_X03_Y0C_lo_unq1),
    .read_config_data(Tile_X03_Y0C_read_config_data),
    .read_config_data_in(Tile_X03_Y0B_read_config_data),
    .reset(Tile_X03_Y0B_reset_out),
    .reset_out(Tile_X03_Y0C_reset_out),
    .stall(Tile_X03_Y0B_stall_out),
    .stall_out(Tile_X03_Y0C_stall_out),
    .tile_id(Tile_X03_Y0C_tile_id_in)
);
mantle_wire__typeBit9 Tile_X03_Y0C_hi (
    .in(Tile_X03_Y0C_hi_unq1),
    .out(Tile_X03_Y0C_hi_out)
);
mantle_wire__typeBit8 Tile_X03_Y0C_lo (
    .in(Tile_X03_Y0C_lo_unq1),
    .out(Tile_X03_Y0C_lo_out)
);
wire [15:0] Tile_X03_Y0C_tile_id_out;
assign Tile_X03_Y0C_tile_id_out = {Tile_X03_Y0C_lo_out[7],Tile_X03_Y0C_lo_out[7:6],Tile_X03_Y0C_lo_out[6:5],Tile_X03_Y0C_lo_out[5],Tile_X03_Y0C_hi_out[5:4],Tile_X03_Y0C_lo_out[3],Tile_X03_Y0C_lo_out[3:2],Tile_X03_Y0C_lo_out[2],Tile_X03_Y0C_hi_out[2:1],Tile_X03_Y0C_lo_out[0],Tile_X03_Y0C_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X03_Y0C_tile_id (
    .in(Tile_X03_Y0C_tile_id_in),
    .out(Tile_X03_Y0C_tile_id_out)
);
Tile_MemCore Tile_X03_Y0D (
    .SB_T0_EAST_SB_IN_B1(Tile_X04_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X04_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X03_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X03_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X03_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X03_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X02_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X02_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X03_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X03_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X04_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X04_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X03_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X03_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X03_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X03_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X02_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X02_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X03_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X03_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X04_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X04_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X03_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X03_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X03_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X03_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X02_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X02_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X03_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X03_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X04_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X04_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X03_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X03_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X03_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X03_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X03_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X03_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X03_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X03_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X02_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X02_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X03_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X03_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X04_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X04_Y0D_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X03_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X03_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X03_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X03_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X03_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X03_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X03_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X03_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X02_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X02_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X03_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X03_Y0D_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y0D_clk_pass_through_out_right),
    .clk_out(Tile_X03_Y0D_clk_out),
    .config_config_addr(Tile_X03_Y0C_config_out_config_addr),
    .config_config_data(Tile_X03_Y0C_config_out_config_data),
    .config_out_config_addr(Tile_X03_Y0D_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y0D_config_out_config_data),
    .config_out_read(Tile_X03_Y0D_config_out_read),
    .config_out_write(Tile_X03_Y0D_config_out_write),
    .config_read(Tile_X03_Y0C_config_out_read),
    .config_write(Tile_X03_Y0C_config_out_write),
    .hi(Tile_X03_Y0D_hi_unq1),
    .lo(Tile_X03_Y0D_lo_unq1),
    .read_config_data(Tile_X03_Y0D_read_config_data),
    .read_config_data_in(Tile_X03_Y0C_read_config_data),
    .reset(Tile_X03_Y0C_reset_out),
    .reset_out(Tile_X03_Y0D_reset_out),
    .stall(Tile_X03_Y0C_stall_out),
    .stall_out(Tile_X03_Y0D_stall_out),
    .tile_id(Tile_X03_Y0D_tile_id_in)
);
mantle_wire__typeBit9 Tile_X03_Y0D_hi (
    .in(Tile_X03_Y0D_hi_unq1),
    .out(Tile_X03_Y0D_hi_out)
);
mantle_wire__typeBit8 Tile_X03_Y0D_lo (
    .in(Tile_X03_Y0D_lo_unq1),
    .out(Tile_X03_Y0D_lo_out)
);
wire [15:0] Tile_X03_Y0D_tile_id_out;
assign Tile_X03_Y0D_tile_id_out = {Tile_X03_Y0D_lo_out[7],Tile_X03_Y0D_lo_out[7:6],Tile_X03_Y0D_lo_out[6:5],Tile_X03_Y0D_lo_out[5],Tile_X03_Y0D_hi_out[5:4],Tile_X03_Y0D_lo_out[3],Tile_X03_Y0D_lo_out[3:2],Tile_X03_Y0D_lo_out[2],Tile_X03_Y0D_hi_out[2:1],Tile_X03_Y0D_lo_out[0],Tile_X03_Y0D_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X03_Y0D_tile_id (
    .in(Tile_X03_Y0D_tile_id_in),
    .out(Tile_X03_Y0D_tile_id_out)
);
Tile_MemCore Tile_X03_Y0E (
    .SB_T0_EAST_SB_IN_B1(Tile_X04_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X04_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X03_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X03_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X03_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X03_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X02_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X02_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X03_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X03_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X04_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X04_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X03_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X03_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X03_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X03_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X02_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X02_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X03_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X03_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X04_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X04_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X03_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X03_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X03_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X03_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X02_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X02_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X03_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X03_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X04_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X04_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X03_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X03_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X03_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X03_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X03_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X03_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X03_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X03_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X02_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X02_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X03_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X03_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X04_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X04_Y0E_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X03_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X03_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X03_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X03_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X03_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X03_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X03_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X03_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X02_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X02_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X03_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X03_Y0E_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y0E_clk_pass_through_out_right),
    .clk_out(Tile_X03_Y0E_clk_out),
    .config_config_addr(Tile_X03_Y0D_config_out_config_addr),
    .config_config_data(Tile_X03_Y0D_config_out_config_data),
    .config_out_config_addr(Tile_X03_Y0E_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y0E_config_out_config_data),
    .config_out_read(Tile_X03_Y0E_config_out_read),
    .config_out_write(Tile_X03_Y0E_config_out_write),
    .config_read(Tile_X03_Y0D_config_out_read),
    .config_write(Tile_X03_Y0D_config_out_write),
    .hi(Tile_X03_Y0E_hi_unq1),
    .lo(Tile_X03_Y0E_lo_unq1),
    .read_config_data(Tile_X03_Y0E_read_config_data),
    .read_config_data_in(Tile_X03_Y0D_read_config_data),
    .reset(Tile_X03_Y0D_reset_out),
    .reset_out(Tile_X03_Y0E_reset_out),
    .stall(Tile_X03_Y0D_stall_out),
    .stall_out(Tile_X03_Y0E_stall_out),
    .tile_id(Tile_X03_Y0E_tile_id_in)
);
mantle_wire__typeBit9 Tile_X03_Y0E_hi (
    .in(Tile_X03_Y0E_hi_unq1),
    .out(Tile_X03_Y0E_hi_out)
);
mantle_wire__typeBit8 Tile_X03_Y0E_lo (
    .in(Tile_X03_Y0E_lo_unq1),
    .out(Tile_X03_Y0E_lo_out)
);
wire [15:0] Tile_X03_Y0E_tile_id_out;
assign Tile_X03_Y0E_tile_id_out = {Tile_X03_Y0E_lo_out[7],Tile_X03_Y0E_lo_out[7:6],Tile_X03_Y0E_lo_out[6:5],Tile_X03_Y0E_lo_out[5],Tile_X03_Y0E_hi_out[5:4],Tile_X03_Y0E_lo_out[3],Tile_X03_Y0E_lo_out[3:2],Tile_X03_Y0E_lo_out[2],Tile_X03_Y0E_hi_out[2:1],Tile_X03_Y0E_hi_out[1],Tile_X03_Y0E_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X03_Y0E_tile_id (
    .in(Tile_X03_Y0E_tile_id_in),
    .out(Tile_X03_Y0E_tile_id_out)
);
Tile_MemCore Tile_X03_Y0F (
    .SB_T0_EAST_SB_IN_B1(Tile_X04_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X04_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X03_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X03_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X03_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X03_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X03_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X03_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X02_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X02_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X03_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X03_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X04_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X04_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X03_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X03_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X03_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X03_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X03_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X03_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X02_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X02_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X03_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X03_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X04_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X04_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X03_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X03_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X03_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X03_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X03_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X03_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X02_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X02_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X03_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X03_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X04_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X04_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X03_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X03_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X03_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X03_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X03_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X03_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X03_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X03_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X02_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X02_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X03_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X03_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X04_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X04_Y0F_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X03_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X03_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X03_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X03_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X03_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X03_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X03_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X03_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X02_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X02_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X03_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X03_Y0F_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y0F_clk_pass_through_out_right),
    .clk_out(Tile_X03_Y0F_clk_out),
    .config_config_addr(Tile_X03_Y0E_config_out_config_addr),
    .config_config_data(Tile_X03_Y0E_config_out_config_data),
    .config_out_config_addr(Tile_X03_Y0F_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y0F_config_out_config_data),
    .config_out_read(Tile_X03_Y0F_config_out_read),
    .config_out_write(Tile_X03_Y0F_config_out_write),
    .config_read(Tile_X03_Y0E_config_out_read),
    .config_write(Tile_X03_Y0E_config_out_write),
    .hi(Tile_X03_Y0F_hi_unq1),
    .lo(Tile_X03_Y0F_lo_unq1),
    .read_config_data(Tile_X03_Y0F_read_config_data),
    .read_config_data_in(Tile_X03_Y0E_read_config_data),
    .reset(Tile_X03_Y0E_reset_out),
    .reset_out(Tile_X03_Y0F_reset_out),
    .stall(Tile_X03_Y0E_stall_out),
    .stall_out(Tile_X03_Y0F_stall_out),
    .tile_id(Tile_X03_Y0F_tile_id_in)
);
mantle_wire__typeBit9 Tile_X03_Y0F_hi (
    .in(Tile_X03_Y0F_hi_unq1),
    .out(Tile_X03_Y0F_hi_out)
);
mantle_wire__typeBit8 Tile_X03_Y0F_lo (
    .in(Tile_X03_Y0F_lo_unq1),
    .out(Tile_X03_Y0F_lo_out)
);
wire [15:0] Tile_X03_Y0F_tile_id_out;
assign Tile_X03_Y0F_tile_id_out = {Tile_X03_Y0F_lo_out[7],Tile_X03_Y0F_lo_out[7:6],Tile_X03_Y0F_lo_out[6:5],Tile_X03_Y0F_lo_out[5],Tile_X03_Y0F_hi_out[5:4],Tile_X03_Y0F_lo_out[3],Tile_X03_Y0F_lo_out[3:2],Tile_X03_Y0F_lo_out[2],Tile_X03_Y0F_hi_out[2:1],Tile_X03_Y0F_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X03_Y0F_tile_id (
    .in(Tile_X03_Y0F_tile_id_in),
    .out(Tile_X03_Y0F_tile_id_out)
);
Tile_MemCore Tile_X03_Y10 (
    .SB_T0_EAST_SB_IN_B1(Tile_X04_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X04_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X03_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X03_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X03_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X03_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X03_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X03_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T0_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X03_Y10_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X03_Y10_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X02_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X02_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X03_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X03_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X04_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X04_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X03_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X03_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X03_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X03_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X03_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X03_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T1_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X03_Y10_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X03_Y10_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X02_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X02_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X03_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X03_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X04_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X04_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X03_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X03_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X03_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X03_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X03_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X03_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T2_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X03_Y10_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X03_Y10_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X02_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X02_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X03_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X03_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X04_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X04_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X03_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X03_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X03_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X03_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X03_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X03_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T3_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X03_Y10_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X03_Y10_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X02_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X02_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X03_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X03_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X04_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X04_Y10_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X03_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X03_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X03_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X03_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X03_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X03_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T4_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X03_Y10_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X03_Y10_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X02_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X02_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X03_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X03_Y10_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X02_Y10_clk_pass_through_out_right),
    .clk_out(Tile_X03_Y10_clk_out),
    .config_config_addr(Tile_X03_Y0F_config_out_config_addr),
    .config_config_data(Tile_X03_Y0F_config_out_config_data),
    .config_out_config_addr(Tile_X03_Y10_config_out_config_addr),
    .config_out_config_data(Tile_X03_Y10_config_out_config_data),
    .config_out_read(Tile_X03_Y10_config_out_read),
    .config_out_write(Tile_X03_Y10_config_out_write),
    .config_read(Tile_X03_Y0F_config_out_read),
    .config_write(Tile_X03_Y0F_config_out_write),
    .hi(Tile_X03_Y10_hi_unq1),
    .lo(Tile_X03_Y10_lo_unq1),
    .read_config_data(Tile_X03_Y10_read_config_data),
    .read_config_data_in(Tile_X03_Y0F_read_config_data),
    .reset(Tile_X03_Y0F_reset_out),
    .reset_out(Tile_X03_Y10_reset_out),
    .stall(Tile_X03_Y0F_stall_out),
    .stall_out(Tile_X03_Y10_stall_out),
    .tile_id(Tile_X03_Y10_tile_id_in)
);
mantle_wire__typeBit9 Tile_X03_Y10_hi (
    .in(Tile_X03_Y10_hi_unq1),
    .out(Tile_X03_Y10_hi_out)
);
mantle_wire__typeBit8 Tile_X03_Y10_lo (
    .in(Tile_X03_Y10_lo_unq1),
    .out(Tile_X03_Y10_lo_out)
);
wire [15:0] Tile_X03_Y10_tile_id_out;
assign Tile_X03_Y10_tile_id_out = {Tile_X03_Y10_lo_out[7],Tile_X03_Y10_lo_out[7:6],Tile_X03_Y10_lo_out[6:5],Tile_X03_Y10_lo_out[5],Tile_X03_Y10_hi_out[5:4],Tile_X03_Y10_lo_out[3],Tile_X03_Y10_lo_out[3:2],Tile_X03_Y10_hi_out[2],Tile_X03_Y10_lo_out[1],Tile_X03_Y10_lo_out[1:0],Tile_X03_Y10_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X03_Y10_tile_id (
    .in(Tile_X03_Y10_tile_id_in),
    .out(Tile_X03_Y10_tile_id_out)
);
wire [15:0] Tile_X04_Y00_tile_id;
assign Tile_X04_Y00_tile_id = {Tile_X04_Y00_lo[7],Tile_X04_Y00_lo[7:6],Tile_X04_Y00_lo[6:5],Tile_X04_Y00_hi[5],Tile_X04_Y00_lo[4],Tile_X04_Y00_lo[4:3],Tile_X04_Y00_lo[3:2],Tile_X04_Y00_lo[2:1],Tile_X04_Y00_lo[1:0],Tile_X04_Y00_lo[0]};
Tile_io_core Tile_X04_Y00 (
    .tile_id(Tile_X04_Y00_tile_id),
    .glb2io_1(glb2io_1_X04_Y00),
    .f2io_1(Tile_X04_Y01_SB_T0_NORTH_SB_OUT_B1),
    .io2glb_1(Tile_X04_Y00_io2glb_1),
    .io2f_1(Tile_X04_Y00_io2f_1),
    .glb2io_16(glb2io_16_X04_Y00),
    .f2io_16(Tile_X04_Y01_SB_T0_NORTH_SB_OUT_B16),
    .io2glb_16(Tile_X04_Y00_io2glb_16),
    .io2f_16(Tile_X04_Y00_io2f_16),
    .hi(Tile_X04_Y00_hi),
    .lo(Tile_X04_Y00_lo)
);
Tile_PE Tile_X04_Y01 (
    .SB_T0_EAST_SB_IN_B1(Tile_X05_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X05_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X04_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X04_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X04_Y00_io2f_1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X04_Y00_io2f_16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X04_Y01_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X04_Y01_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X04_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X04_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X04_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X04_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X03_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X03_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X04_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X04_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X05_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X05_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X04_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X04_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X04_Y00_io2f_1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X04_Y00_io2f_16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X04_Y01_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X04_Y01_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X04_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X04_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X04_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X04_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X03_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X03_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X04_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X04_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X05_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X05_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X04_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X04_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X04_Y00_io2f_1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X04_Y00_io2f_16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X04_Y01_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X04_Y01_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X04_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X04_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X04_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X04_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X03_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X03_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X04_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X04_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X05_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X05_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X04_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X04_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X04_Y00_io2f_1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X04_Y00_io2f_16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X04_Y01_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X04_Y01_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X04_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X04_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X04_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X04_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X03_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X03_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X04_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X04_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X05_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X05_Y01_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X04_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X04_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X04_Y00_io2f_1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X04_Y00_io2f_16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X04_Y01_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X04_Y01_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X04_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X04_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X04_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X04_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X03_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X03_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X04_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X04_Y01_SB_T4_WEST_SB_OUT_B16),
    .clk(clk),
    .clk_out(Tile_X04_Y01_clk_out),
    .clk_pass_through(clk),
    .clk_pass_through_out_bot(Tile_X04_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X04_Y01_clk_pass_through_out_right),
    .config_config_addr(config_4_config_addr),
    .config_config_data(config_4_config_data),
    .config_out_config_addr(Tile_X04_Y01_config_out_config_addr),
    .config_out_config_data(Tile_X04_Y01_config_out_config_data),
    .config_out_read(Tile_X04_Y01_config_out_read),
    .config_out_write(Tile_X04_Y01_config_out_write),
    .config_read(config_4_read),
    .config_write(config_4_write),
    .hi(Tile_X04_Y01_hi),
    .lo(Tile_X04_Y01_lo_unq1),
    .read_config_data(Tile_X04_Y01_read_config_data),
    .read_config_data_in(const_0_32_out),
    .reset(reset),
    .reset_out(Tile_X04_Y01_reset_out),
    .stall(stall[4]),
    .stall_out(Tile_X04_Y01_stall_out),
    .tile_id(Tile_X04_Y01_tile_id_in)
);
mantle_wire__typeBit8 Tile_X04_Y01_lo (
    .in(Tile_X04_Y01_lo_unq1),
    .out(Tile_X04_Y01_lo_out)
);
wire [15:0] Tile_X04_Y01_tile_id_out;
assign Tile_X04_Y01_tile_id_out = {Tile_X04_Y01_lo_out[7],Tile_X04_Y01_lo_out[7:6],Tile_X04_Y01_lo_out[6:5],Tile_X04_Y01_hi[5],Tile_X04_Y01_lo_out[4],Tile_X04_Y01_lo_out[4:3],Tile_X04_Y01_lo_out[3:2],Tile_X04_Y01_lo_out[2:1],Tile_X04_Y01_lo_out[1:0],Tile_X04_Y01_hi[0]};
mantle_wire__typeBitIn16 Tile_X04_Y01_tile_id (
    .in(Tile_X04_Y01_tile_id_in),
    .out(Tile_X04_Y01_tile_id_out)
);
Tile_PE Tile_X04_Y02 (
    .SB_T0_EAST_SB_IN_B1(Tile_X05_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X05_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X04_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X04_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X04_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X04_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X04_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X04_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X04_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X04_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X04_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X04_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X03_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X03_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X04_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X04_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X05_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X05_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X04_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X04_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X04_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X04_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X04_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X04_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X04_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X04_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X04_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X04_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X03_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X03_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X04_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X04_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X05_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X05_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X04_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X04_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X04_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X04_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X04_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X04_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X04_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X04_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X04_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X04_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X03_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X03_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X04_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X04_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X05_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X05_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X04_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X04_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X04_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X04_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X04_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X04_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X04_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X04_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X04_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X04_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X03_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X03_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X04_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X04_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X05_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X05_Y02_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X04_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X04_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X04_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X04_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X04_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X04_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X04_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X04_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X04_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X04_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X03_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X03_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X04_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X04_Y02_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X04_Y01_clk_out),
    .clk_out(Tile_X04_Y02_clk_out),
    .clk_pass_through(Tile_X04_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X04_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X04_Y02_clk_pass_through_out_right),
    .config_config_addr(Tile_X04_Y01_config_out_config_addr),
    .config_config_data(Tile_X04_Y01_config_out_config_data),
    .config_out_config_addr(Tile_X04_Y02_config_out_config_addr),
    .config_out_config_data(Tile_X04_Y02_config_out_config_data),
    .config_out_read(Tile_X04_Y02_config_out_read),
    .config_out_write(Tile_X04_Y02_config_out_write),
    .config_read(Tile_X04_Y01_config_out_read),
    .config_write(Tile_X04_Y01_config_out_write),
    .hi(Tile_X04_Y02_hi),
    .lo(Tile_X04_Y02_lo_unq1),
    .read_config_data(Tile_X04_Y02_read_config_data),
    .read_config_data_in(Tile_X04_Y01_read_config_data),
    .reset(Tile_X04_Y01_reset_out),
    .reset_out(Tile_X04_Y02_reset_out),
    .stall(Tile_X04_Y01_stall_out),
    .stall_out(Tile_X04_Y02_stall_out),
    .tile_id(Tile_X04_Y02_tile_id_in)
);
mantle_wire__typeBit8 Tile_X04_Y02_lo (
    .in(Tile_X04_Y02_lo_unq1),
    .out(Tile_X04_Y02_lo_out)
);
wire [15:0] Tile_X04_Y02_tile_id_out;
assign Tile_X04_Y02_tile_id_out = {Tile_X04_Y02_lo_out[7],Tile_X04_Y02_lo_out[7:6],Tile_X04_Y02_lo_out[6:5],Tile_X04_Y02_hi[5],Tile_X04_Y02_lo_out[4],Tile_X04_Y02_lo_out[4:3],Tile_X04_Y02_lo_out[3:2],Tile_X04_Y02_lo_out[2:1],Tile_X04_Y02_lo_out[1],Tile_X04_Y02_hi[1],Tile_X04_Y02_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X04_Y02_tile_id (
    .in(Tile_X04_Y02_tile_id_in),
    .out(Tile_X04_Y02_tile_id_out)
);
Tile_PE Tile_X04_Y03 (
    .SB_T0_EAST_SB_IN_B1(Tile_X05_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X05_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X04_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X04_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X04_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X04_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X04_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X04_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X04_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X04_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X04_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X04_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X03_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X03_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X04_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X04_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X05_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X05_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X04_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X04_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X04_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X04_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X04_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X04_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X04_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X04_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X04_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X04_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X03_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X03_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X04_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X04_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X05_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X05_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X04_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X04_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X04_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X04_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X04_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X04_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X04_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X04_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X04_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X04_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X03_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X03_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X04_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X04_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X05_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X05_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X04_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X04_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X04_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X04_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X04_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X04_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X04_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X04_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X04_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X04_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X03_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X03_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X04_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X04_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X05_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X05_Y03_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X04_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X04_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X04_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X04_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X04_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X04_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X04_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X04_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X04_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X04_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X03_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X03_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X04_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X04_Y03_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X04_Y02_clk_out),
    .clk_out(Tile_X04_Y03_clk_out),
    .clk_pass_through(Tile_X04_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X04_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X04_Y03_clk_pass_through_out_right),
    .config_config_addr(Tile_X04_Y02_config_out_config_addr),
    .config_config_data(Tile_X04_Y02_config_out_config_data),
    .config_out_config_addr(Tile_X04_Y03_config_out_config_addr),
    .config_out_config_data(Tile_X04_Y03_config_out_config_data),
    .config_out_read(Tile_X04_Y03_config_out_read),
    .config_out_write(Tile_X04_Y03_config_out_write),
    .config_read(Tile_X04_Y02_config_out_read),
    .config_write(Tile_X04_Y02_config_out_write),
    .hi(Tile_X04_Y03_hi_unq1),
    .lo(Tile_X04_Y03_lo_unq1),
    .read_config_data(Tile_X04_Y03_read_config_data),
    .read_config_data_in(Tile_X04_Y02_read_config_data),
    .reset(Tile_X04_Y02_reset_out),
    .reset_out(Tile_X04_Y03_reset_out),
    .stall(Tile_X04_Y02_stall_out),
    .stall_out(Tile_X04_Y03_stall_out),
    .tile_id(Tile_X04_Y03_tile_id_in)
);
mantle_wire__typeBit9 Tile_X04_Y03_hi (
    .in(Tile_X04_Y03_hi_unq1),
    .out(Tile_X04_Y03_hi_out)
);
mantle_wire__typeBit8 Tile_X04_Y03_lo (
    .in(Tile_X04_Y03_lo_unq1),
    .out(Tile_X04_Y03_lo_out)
);
wire [15:0] Tile_X04_Y03_tile_id_out;
assign Tile_X04_Y03_tile_id_out = {Tile_X04_Y03_lo_out[7],Tile_X04_Y03_lo_out[7:6],Tile_X04_Y03_lo_out[6:5],Tile_X04_Y03_hi_out[5],Tile_X04_Y03_lo_out[4],Tile_X04_Y03_lo_out[4:3],Tile_X04_Y03_lo_out[3:2],Tile_X04_Y03_lo_out[2:1],Tile_X04_Y03_lo_out[1],Tile_X04_Y03_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X04_Y03_tile_id (
    .in(Tile_X04_Y03_tile_id_in),
    .out(Tile_X04_Y03_tile_id_out)
);
Tile_PE Tile_X04_Y04 (
    .SB_T0_EAST_SB_IN_B1(Tile_X05_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X05_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X04_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X04_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X04_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X04_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X04_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X04_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X04_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X04_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X04_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X04_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X03_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X03_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X04_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X04_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X05_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X05_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X04_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X04_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X04_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X04_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X04_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X04_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X04_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X04_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X04_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X04_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X03_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X03_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X04_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X04_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X05_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X05_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X04_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X04_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X04_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X04_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X04_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X04_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X04_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X04_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X04_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X04_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X03_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X03_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X04_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X04_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X05_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X05_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X04_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X04_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X04_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X04_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X04_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X04_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X04_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X04_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X04_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X04_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X03_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X03_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X04_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X04_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X05_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X05_Y04_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X04_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X04_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X04_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X04_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X04_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X04_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X04_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X04_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X04_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X04_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X03_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X03_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X04_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X04_Y04_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X04_Y03_clk_out),
    .clk_out(Tile_X04_Y04_clk_out),
    .clk_pass_through(Tile_X04_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X04_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X04_Y04_clk_pass_through_out_right),
    .config_config_addr(Tile_X04_Y03_config_out_config_addr),
    .config_config_data(Tile_X04_Y03_config_out_config_data),
    .config_out_config_addr(Tile_X04_Y04_config_out_config_addr),
    .config_out_config_data(Tile_X04_Y04_config_out_config_data),
    .config_out_read(Tile_X04_Y04_config_out_read),
    .config_out_write(Tile_X04_Y04_config_out_write),
    .config_read(Tile_X04_Y03_config_out_read),
    .config_write(Tile_X04_Y03_config_out_write),
    .hi(Tile_X04_Y04_hi),
    .lo(Tile_X04_Y04_lo_unq1),
    .read_config_data(Tile_X04_Y04_read_config_data),
    .read_config_data_in(Tile_X04_Y03_read_config_data),
    .reset(Tile_X04_Y03_reset_out),
    .reset_out(Tile_X04_Y04_reset_out),
    .stall(Tile_X04_Y03_stall_out),
    .stall_out(Tile_X04_Y04_stall_out),
    .tile_id(Tile_X04_Y04_tile_id_in)
);
mantle_wire__typeBit8 Tile_X04_Y04_lo (
    .in(Tile_X04_Y04_lo_unq1),
    .out(Tile_X04_Y04_lo_out)
);
wire [15:0] Tile_X04_Y04_tile_id_out;
assign Tile_X04_Y04_tile_id_out = {Tile_X04_Y04_lo_out[7],Tile_X04_Y04_lo_out[7:6],Tile_X04_Y04_lo_out[6:5],Tile_X04_Y04_hi[5],Tile_X04_Y04_lo_out[4],Tile_X04_Y04_lo_out[4:3],Tile_X04_Y04_lo_out[3:2],Tile_X04_Y04_lo_out[2:1],Tile_X04_Y04_hi[1],Tile_X04_Y04_lo_out[0],Tile_X04_Y04_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X04_Y04_tile_id (
    .in(Tile_X04_Y04_tile_id_in),
    .out(Tile_X04_Y04_tile_id_out)
);
Tile_PE Tile_X04_Y05 (
    .SB_T0_EAST_SB_IN_B1(Tile_X05_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X05_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X04_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X04_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X04_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X04_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X04_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X04_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X04_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X04_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X04_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X04_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X03_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X03_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X04_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X04_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X05_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X05_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X04_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X04_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X04_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X04_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X04_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X04_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X04_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X04_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X04_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X04_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X03_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X03_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X04_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X04_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X05_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X05_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X04_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X04_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X04_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X04_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X04_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X04_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X04_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X04_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X04_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X04_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X03_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X03_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X04_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X04_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X05_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X05_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X04_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X04_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X04_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X04_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X04_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X04_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X04_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X04_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X04_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X04_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X03_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X03_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X04_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X04_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X05_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X05_Y05_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X04_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X04_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X04_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X04_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X04_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X04_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X04_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X04_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X04_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X04_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X03_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X03_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X04_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X04_Y05_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X04_Y04_clk_out),
    .clk_out(Tile_X04_Y05_clk_out),
    .clk_pass_through(Tile_X04_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X04_Y05_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X04_Y05_clk_pass_through_out_right),
    .config_config_addr(Tile_X04_Y04_config_out_config_addr),
    .config_config_data(Tile_X04_Y04_config_out_config_data),
    .config_out_config_addr(Tile_X04_Y05_config_out_config_addr),
    .config_out_config_data(Tile_X04_Y05_config_out_config_data),
    .config_out_read(Tile_X04_Y05_config_out_read),
    .config_out_write(Tile_X04_Y05_config_out_write),
    .config_read(Tile_X04_Y04_config_out_read),
    .config_write(Tile_X04_Y04_config_out_write),
    .hi(Tile_X04_Y05_hi),
    .lo(Tile_X04_Y05_lo_unq1),
    .read_config_data(Tile_X04_Y05_read_config_data),
    .read_config_data_in(Tile_X04_Y04_read_config_data),
    .reset(Tile_X04_Y04_reset_out),
    .reset_out(Tile_X04_Y05_reset_out),
    .stall(Tile_X04_Y04_stall_out),
    .stall_out(Tile_X04_Y05_stall_out),
    .tile_id(Tile_X04_Y05_tile_id_in)
);
mantle_wire__typeBit8 Tile_X04_Y05_lo (
    .in(Tile_X04_Y05_lo_unq1),
    .out(Tile_X04_Y05_lo_out)
);
wire [15:0] Tile_X04_Y05_tile_id_out;
assign Tile_X04_Y05_tile_id_out = {Tile_X04_Y05_lo_out[7],Tile_X04_Y05_lo_out[7:6],Tile_X04_Y05_lo_out[6:5],Tile_X04_Y05_hi[5],Tile_X04_Y05_lo_out[4],Tile_X04_Y05_lo_out[4:3],Tile_X04_Y05_lo_out[3:2],Tile_X04_Y05_lo_out[2:1],Tile_X04_Y05_hi[1],Tile_X04_Y05_lo_out[0],Tile_X04_Y05_hi[0]};
mantle_wire__typeBitIn16 Tile_X04_Y05_tile_id (
    .in(Tile_X04_Y05_tile_id_in),
    .out(Tile_X04_Y05_tile_id_out)
);
Tile_PE Tile_X04_Y06 (
    .SB_T0_EAST_SB_IN_B1(Tile_X05_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X05_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X04_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X04_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X04_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X04_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X04_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X04_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X04_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X04_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X04_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X04_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X03_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X03_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X04_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X04_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X05_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X05_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X04_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X04_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X04_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X04_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X04_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X04_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X04_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X04_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X04_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X04_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X03_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X03_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X04_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X04_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X05_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X05_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X04_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X04_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X04_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X04_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X04_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X04_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X04_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X04_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X04_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X04_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X03_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X03_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X04_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X04_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X05_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X05_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X04_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X04_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X04_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X04_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X04_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X04_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X04_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X04_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X04_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X04_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X03_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X03_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X04_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X04_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X05_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X05_Y06_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X04_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X04_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X04_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X04_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X04_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X04_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X04_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X04_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X04_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X04_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X03_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X03_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X04_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X04_Y06_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X04_Y05_clk_out),
    .clk_out(Tile_X04_Y06_clk_out),
    .clk_pass_through(Tile_X04_Y05_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X04_Y06_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X04_Y06_clk_pass_through_out_right),
    .config_config_addr(Tile_X04_Y05_config_out_config_addr),
    .config_config_data(Tile_X04_Y05_config_out_config_data),
    .config_out_config_addr(Tile_X04_Y06_config_out_config_addr),
    .config_out_config_data(Tile_X04_Y06_config_out_config_data),
    .config_out_read(Tile_X04_Y06_config_out_read),
    .config_out_write(Tile_X04_Y06_config_out_write),
    .config_read(Tile_X04_Y05_config_out_read),
    .config_write(Tile_X04_Y05_config_out_write),
    .hi(Tile_X04_Y06_hi),
    .lo(Tile_X04_Y06_lo_unq1),
    .read_config_data(Tile_X04_Y06_read_config_data),
    .read_config_data_in(Tile_X04_Y05_read_config_data),
    .reset(Tile_X04_Y05_reset_out),
    .reset_out(Tile_X04_Y06_reset_out),
    .stall(Tile_X04_Y05_stall_out),
    .stall_out(Tile_X04_Y06_stall_out),
    .tile_id(Tile_X04_Y06_tile_id_in)
);
mantle_wire__typeBit8 Tile_X04_Y06_lo (
    .in(Tile_X04_Y06_lo_unq1),
    .out(Tile_X04_Y06_lo_out)
);
wire [15:0] Tile_X04_Y06_tile_id_out;
assign Tile_X04_Y06_tile_id_out = {Tile_X04_Y06_lo_out[7],Tile_X04_Y06_lo_out[7:6],Tile_X04_Y06_lo_out[6:5],Tile_X04_Y06_hi[5],Tile_X04_Y06_lo_out[4],Tile_X04_Y06_lo_out[4:3],Tile_X04_Y06_lo_out[3:2],Tile_X04_Y06_lo_out[2:1],Tile_X04_Y06_hi[1],Tile_X04_Y06_hi[1],Tile_X04_Y06_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X04_Y06_tile_id (
    .in(Tile_X04_Y06_tile_id_in),
    .out(Tile_X04_Y06_tile_id_out)
);
Tile_PE Tile_X04_Y07 (
    .SB_T0_EAST_SB_IN_B1(Tile_X05_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X05_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X04_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X04_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X04_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X04_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X04_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X04_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X04_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X04_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X04_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X04_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X03_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X03_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X04_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X04_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X05_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X05_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X04_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X04_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X04_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X04_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X04_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X04_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X04_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X04_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X04_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X04_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X03_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X03_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X04_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X04_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X05_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X05_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X04_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X04_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X04_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X04_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X04_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X04_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X04_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X04_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X04_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X04_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X03_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X03_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X04_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X04_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X05_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X05_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X04_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X04_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X04_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X04_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X04_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X04_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X04_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X04_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X04_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X04_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X03_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X03_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X04_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X04_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X05_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X05_Y07_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X04_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X04_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X04_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X04_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X04_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X04_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X04_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X04_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X04_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X04_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X03_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X03_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X04_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X04_Y07_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X04_Y06_clk_out),
    .clk_out(Tile_X04_Y07_clk_out),
    .clk_pass_through(Tile_X04_Y06_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X04_Y07_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X04_Y07_clk_pass_through_out_right),
    .config_config_addr(Tile_X04_Y06_config_out_config_addr),
    .config_config_data(Tile_X04_Y06_config_out_config_data),
    .config_out_config_addr(Tile_X04_Y07_config_out_config_addr),
    .config_out_config_data(Tile_X04_Y07_config_out_config_data),
    .config_out_read(Tile_X04_Y07_config_out_read),
    .config_out_write(Tile_X04_Y07_config_out_write),
    .config_read(Tile_X04_Y06_config_out_read),
    .config_write(Tile_X04_Y06_config_out_write),
    .hi(Tile_X04_Y07_hi_unq1),
    .lo(Tile_X04_Y07_lo_unq1),
    .read_config_data(Tile_X04_Y07_read_config_data),
    .read_config_data_in(Tile_X04_Y06_read_config_data),
    .reset(Tile_X04_Y06_reset_out),
    .reset_out(Tile_X04_Y07_reset_out),
    .stall(Tile_X04_Y06_stall_out),
    .stall_out(Tile_X04_Y07_stall_out),
    .tile_id(Tile_X04_Y07_tile_id_in)
);
mantle_wire__typeBit9 Tile_X04_Y07_hi (
    .in(Tile_X04_Y07_hi_unq1),
    .out(Tile_X04_Y07_hi_out)
);
mantle_wire__typeBit8 Tile_X04_Y07_lo (
    .in(Tile_X04_Y07_lo_unq1),
    .out(Tile_X04_Y07_lo_out)
);
wire [15:0] Tile_X04_Y07_tile_id_out;
assign Tile_X04_Y07_tile_id_out = {Tile_X04_Y07_lo_out[7],Tile_X04_Y07_lo_out[7:6],Tile_X04_Y07_lo_out[6:5],Tile_X04_Y07_hi_out[5],Tile_X04_Y07_lo_out[4],Tile_X04_Y07_lo_out[4:3],Tile_X04_Y07_lo_out[3:2],Tile_X04_Y07_lo_out[2:1],Tile_X04_Y07_hi_out[1],Tile_X04_Y07_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X04_Y07_tile_id (
    .in(Tile_X04_Y07_tile_id_in),
    .out(Tile_X04_Y07_tile_id_out)
);
Tile_PE Tile_X04_Y08 (
    .SB_T0_EAST_SB_IN_B1(Tile_X05_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X05_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X04_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X04_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X04_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X04_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X04_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X04_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X04_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X04_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X04_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X04_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X03_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X03_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X04_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X04_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X05_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X05_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X04_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X04_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X04_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X04_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X04_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X04_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X04_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X04_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X04_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X04_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X03_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X03_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X04_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X04_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X05_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X05_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X04_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X04_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X04_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X04_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X04_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X04_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X04_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X04_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X04_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X04_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X03_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X03_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X04_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X04_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X05_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X05_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X04_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X04_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X04_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X04_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X04_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X04_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X04_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X04_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X04_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X04_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X03_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X03_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X04_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X04_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X05_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X05_Y08_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X04_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X04_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X04_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X04_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X04_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X04_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X04_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X04_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X04_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X04_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X03_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X03_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X04_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X04_Y08_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X04_Y07_clk_out),
    .clk_out(Tile_X04_Y08_clk_out),
    .clk_pass_through(Tile_X04_Y07_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X04_Y08_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X04_Y08_clk_pass_through_out_right),
    .config_config_addr(Tile_X04_Y07_config_out_config_addr),
    .config_config_data(Tile_X04_Y07_config_out_config_data),
    .config_out_config_addr(Tile_X04_Y08_config_out_config_addr),
    .config_out_config_data(Tile_X04_Y08_config_out_config_data),
    .config_out_read(Tile_X04_Y08_config_out_read),
    .config_out_write(Tile_X04_Y08_config_out_write),
    .config_read(Tile_X04_Y07_config_out_read),
    .config_write(Tile_X04_Y07_config_out_write),
    .hi(Tile_X04_Y08_hi),
    .lo(Tile_X04_Y08_lo_unq1),
    .read_config_data(Tile_X04_Y08_read_config_data),
    .read_config_data_in(Tile_X04_Y07_read_config_data),
    .reset(Tile_X04_Y07_reset_out),
    .reset_out(Tile_X04_Y08_reset_out),
    .stall(Tile_X04_Y07_stall_out),
    .stall_out(Tile_X04_Y08_stall_out),
    .tile_id(Tile_X04_Y08_tile_id_in)
);
mantle_wire__typeBit8 Tile_X04_Y08_lo (
    .in(Tile_X04_Y08_lo_unq1),
    .out(Tile_X04_Y08_lo_out)
);
wire [15:0] Tile_X04_Y08_tile_id_out;
assign Tile_X04_Y08_tile_id_out = {Tile_X04_Y08_lo_out[7],Tile_X04_Y08_lo_out[7:6],Tile_X04_Y08_lo_out[6:5],Tile_X04_Y08_hi[5],Tile_X04_Y08_lo_out[4],Tile_X04_Y08_lo_out[4:3],Tile_X04_Y08_lo_out[3:2],Tile_X04_Y08_lo_out[2],Tile_X04_Y08_hi[2],Tile_X04_Y08_lo_out[1:0],Tile_X04_Y08_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X04_Y08_tile_id (
    .in(Tile_X04_Y08_tile_id_in),
    .out(Tile_X04_Y08_tile_id_out)
);
Tile_PE Tile_X04_Y09 (
    .SB_T0_EAST_SB_IN_B1(Tile_X05_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X05_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X04_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X04_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X04_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X04_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X04_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X04_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X04_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X04_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X04_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X04_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X03_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X03_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X04_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X04_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X05_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X05_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X04_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X04_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X04_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X04_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X04_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X04_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X04_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X04_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X04_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X04_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X03_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X03_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X04_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X04_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X05_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X05_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X04_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X04_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X04_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X04_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X04_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X04_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X04_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X04_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X04_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X04_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X03_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X03_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X04_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X04_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X05_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X05_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X04_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X04_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X04_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X04_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X04_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X04_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X04_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X04_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X04_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X04_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X03_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X03_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X04_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X04_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X05_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X05_Y09_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X04_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X04_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X04_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X04_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X04_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X04_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X04_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X04_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X04_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X04_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X03_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X03_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X04_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X04_Y09_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X04_Y08_clk_out),
    .clk_out(Tile_X04_Y09_clk_out),
    .clk_pass_through(Tile_X04_Y08_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X04_Y09_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X04_Y09_clk_pass_through_out_right),
    .config_config_addr(ConfigPipeStage_inst4_config_out_config_addr),
    .config_config_data(ConfigPipeStage_inst4_config_out_config_data),
    .config_out_config_addr(Tile_X04_Y09_config_out_config_addr),
    .config_out_config_data(Tile_X04_Y09_config_out_config_data),
    .config_out_read(Tile_X04_Y09_config_out_read),
    .config_out_write(Tile_X04_Y09_config_out_write),
    .config_read(ConfigPipeStage_inst4_config_out_read),
    .config_write(ConfigPipeStage_inst4_config_out_write),
    .hi(Tile_X04_Y09_hi),
    .lo(Tile_X04_Y09_lo_unq1),
    .read_config_data(Tile_X04_Y09_read_config_data),
    .read_config_data_in(Tile_X04_Y08_read_config_data),
    .reset(Tile_X04_Y08_reset_out),
    .reset_out(Tile_X04_Y09_reset_out),
    .stall(Tile_X04_Y08_stall_out),
    .stall_out(Tile_X04_Y09_stall_out),
    .tile_id(Tile_X04_Y09_tile_id_in)
);
mantle_wire__typeBit8 Tile_X04_Y09_lo (
    .in(Tile_X04_Y09_lo_unq1),
    .out(Tile_X04_Y09_lo_out)
);
wire [15:0] Tile_X04_Y09_tile_id_out;
assign Tile_X04_Y09_tile_id_out = {Tile_X04_Y09_lo_out[7],Tile_X04_Y09_lo_out[7:6],Tile_X04_Y09_lo_out[6:5],Tile_X04_Y09_hi[5],Tile_X04_Y09_lo_out[4],Tile_X04_Y09_lo_out[4:3],Tile_X04_Y09_lo_out[3:2],Tile_X04_Y09_lo_out[2],Tile_X04_Y09_hi[2],Tile_X04_Y09_lo_out[1:0],Tile_X04_Y09_hi[0]};
mantle_wire__typeBitIn16 Tile_X04_Y09_tile_id (
    .in(Tile_X04_Y09_tile_id_in),
    .out(Tile_X04_Y09_tile_id_out)
);
Tile_PE Tile_X04_Y0A (
    .SB_T0_EAST_SB_IN_B1(Tile_X05_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X05_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X04_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X04_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X04_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X04_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X04_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X04_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X04_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X04_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X04_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X04_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X03_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X03_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X04_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X04_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X05_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X05_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X04_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X04_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X04_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X04_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X04_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X04_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X04_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X04_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X04_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X04_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X03_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X03_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X04_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X04_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X05_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X05_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X04_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X04_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X04_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X04_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X04_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X04_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X04_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X04_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X04_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X04_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X03_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X03_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X04_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X04_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X05_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X05_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X04_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X04_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X04_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X04_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X04_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X04_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X04_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X04_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X04_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X04_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X03_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X03_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X04_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X04_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X05_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X05_Y0A_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X04_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X04_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X04_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X04_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X04_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X04_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X04_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X04_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X04_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X04_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X03_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X03_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X04_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X04_Y0A_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X04_Y09_clk_out),
    .clk_out(Tile_X04_Y0A_clk_out),
    .clk_pass_through(Tile_X04_Y09_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X04_Y0A_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X04_Y0A_clk_pass_through_out_right),
    .config_config_addr(Tile_X04_Y09_config_out_config_addr),
    .config_config_data(Tile_X04_Y09_config_out_config_data),
    .config_out_config_addr(Tile_X04_Y0A_config_out_config_addr),
    .config_out_config_data(Tile_X04_Y0A_config_out_config_data),
    .config_out_read(Tile_X04_Y0A_config_out_read),
    .config_out_write(Tile_X04_Y0A_config_out_write),
    .config_read(Tile_X04_Y09_config_out_read),
    .config_write(Tile_X04_Y09_config_out_write),
    .hi(Tile_X04_Y0A_hi),
    .lo(Tile_X04_Y0A_lo_unq1),
    .read_config_data(Tile_X04_Y0A_read_config_data),
    .read_config_data_in(Tile_X04_Y09_read_config_data),
    .reset(Tile_X04_Y09_reset_out),
    .reset_out(Tile_X04_Y0A_reset_out),
    .stall(Tile_X04_Y09_stall_out),
    .stall_out(Tile_X04_Y0A_stall_out),
    .tile_id(Tile_X04_Y0A_tile_id_in)
);
mantle_wire__typeBit8 Tile_X04_Y0A_lo (
    .in(Tile_X04_Y0A_lo_unq1),
    .out(Tile_X04_Y0A_lo_out)
);
wire [15:0] Tile_X04_Y0A_tile_id_out;
assign Tile_X04_Y0A_tile_id_out = {Tile_X04_Y0A_lo_out[7],Tile_X04_Y0A_lo_out[7:6],Tile_X04_Y0A_lo_out[6:5],Tile_X04_Y0A_hi[5],Tile_X04_Y0A_lo_out[4],Tile_X04_Y0A_lo_out[4:3],Tile_X04_Y0A_lo_out[3:2],Tile_X04_Y0A_lo_out[2],Tile_X04_Y0A_hi[2],Tile_X04_Y0A_lo_out[1],Tile_X04_Y0A_hi[1],Tile_X04_Y0A_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X04_Y0A_tile_id (
    .in(Tile_X04_Y0A_tile_id_in),
    .out(Tile_X04_Y0A_tile_id_out)
);
Tile_PE Tile_X04_Y0B (
    .SB_T0_EAST_SB_IN_B1(Tile_X05_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X05_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X04_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X04_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X04_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X04_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X04_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X04_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X04_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X04_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X04_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X04_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X03_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X03_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X04_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X04_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X05_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X05_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X04_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X04_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X04_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X04_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X04_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X04_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X04_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X04_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X04_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X04_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X03_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X03_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X04_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X04_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X05_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X05_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X04_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X04_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X04_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X04_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X04_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X04_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X04_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X04_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X04_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X04_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X03_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X03_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X04_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X04_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X05_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X05_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X04_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X04_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X04_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X04_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X04_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X04_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X04_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X04_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X04_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X04_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X03_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X03_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X04_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X04_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X05_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X05_Y0B_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X04_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X04_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X04_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X04_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X04_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X04_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X04_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X04_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X04_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X04_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X03_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X03_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X04_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X04_Y0B_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X04_Y0A_clk_out),
    .clk_out(Tile_X04_Y0B_clk_out),
    .clk_pass_through(Tile_X04_Y0A_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X04_Y0B_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X04_Y0B_clk_pass_through_out_right),
    .config_config_addr(Tile_X04_Y0A_config_out_config_addr),
    .config_config_data(Tile_X04_Y0A_config_out_config_data),
    .config_out_config_addr(Tile_X04_Y0B_config_out_config_addr),
    .config_out_config_data(Tile_X04_Y0B_config_out_config_data),
    .config_out_read(Tile_X04_Y0B_config_out_read),
    .config_out_write(Tile_X04_Y0B_config_out_write),
    .config_read(Tile_X04_Y0A_config_out_read),
    .config_write(Tile_X04_Y0A_config_out_write),
    .hi(Tile_X04_Y0B_hi_unq1),
    .lo(Tile_X04_Y0B_lo_unq1),
    .read_config_data(Tile_X04_Y0B_read_config_data),
    .read_config_data_in(Tile_X04_Y0A_read_config_data),
    .reset(Tile_X04_Y0A_reset_out),
    .reset_out(Tile_X04_Y0B_reset_out),
    .stall(Tile_X04_Y0A_stall_out),
    .stall_out(Tile_X04_Y0B_stall_out),
    .tile_id(Tile_X04_Y0B_tile_id_in)
);
mantle_wire__typeBit9 Tile_X04_Y0B_hi (
    .in(Tile_X04_Y0B_hi_unq1),
    .out(Tile_X04_Y0B_hi_out)
);
mantle_wire__typeBit8 Tile_X04_Y0B_lo (
    .in(Tile_X04_Y0B_lo_unq1),
    .out(Tile_X04_Y0B_lo_out)
);
wire [15:0] Tile_X04_Y0B_tile_id_out;
assign Tile_X04_Y0B_tile_id_out = {Tile_X04_Y0B_lo_out[7],Tile_X04_Y0B_lo_out[7:6],Tile_X04_Y0B_lo_out[6:5],Tile_X04_Y0B_hi_out[5],Tile_X04_Y0B_lo_out[4],Tile_X04_Y0B_lo_out[4:3],Tile_X04_Y0B_lo_out[3:2],Tile_X04_Y0B_lo_out[2],Tile_X04_Y0B_hi_out[2],Tile_X04_Y0B_lo_out[1],Tile_X04_Y0B_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X04_Y0B_tile_id (
    .in(Tile_X04_Y0B_tile_id_in),
    .out(Tile_X04_Y0B_tile_id_out)
);
Tile_PE Tile_X04_Y0C (
    .SB_T0_EAST_SB_IN_B1(Tile_X05_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X05_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X04_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X04_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X04_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X04_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X04_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X04_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X04_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X04_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X04_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X04_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X03_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X03_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X04_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X04_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X05_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X05_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X04_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X04_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X04_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X04_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X04_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X04_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X04_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X04_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X04_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X04_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X03_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X03_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X04_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X04_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X05_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X05_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X04_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X04_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X04_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X04_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X04_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X04_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X04_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X04_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X04_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X04_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X03_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X03_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X04_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X04_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X05_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X05_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X04_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X04_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X04_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X04_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X04_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X04_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X04_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X04_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X04_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X04_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X03_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X03_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X04_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X04_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X05_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X05_Y0C_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X04_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X04_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X04_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X04_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X04_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X04_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X04_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X04_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X04_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X04_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X03_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X03_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X04_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X04_Y0C_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X04_Y0B_clk_out),
    .clk_out(Tile_X04_Y0C_clk_out),
    .clk_pass_through(Tile_X04_Y0B_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X04_Y0C_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X04_Y0C_clk_pass_through_out_right),
    .config_config_addr(Tile_X04_Y0B_config_out_config_addr),
    .config_config_data(Tile_X04_Y0B_config_out_config_data),
    .config_out_config_addr(Tile_X04_Y0C_config_out_config_addr),
    .config_out_config_data(Tile_X04_Y0C_config_out_config_data),
    .config_out_read(Tile_X04_Y0C_config_out_read),
    .config_out_write(Tile_X04_Y0C_config_out_write),
    .config_read(Tile_X04_Y0B_config_out_read),
    .config_write(Tile_X04_Y0B_config_out_write),
    .hi(Tile_X04_Y0C_hi_unq1),
    .lo(Tile_X04_Y0C_lo_unq1),
    .read_config_data(Tile_X04_Y0C_read_config_data),
    .read_config_data_in(Tile_X04_Y0B_read_config_data),
    .reset(Tile_X04_Y0B_reset_out),
    .reset_out(Tile_X04_Y0C_reset_out),
    .stall(Tile_X04_Y0B_stall_out),
    .stall_out(Tile_X04_Y0C_stall_out),
    .tile_id(Tile_X04_Y0C_tile_id_in)
);
mantle_wire__typeBit9 Tile_X04_Y0C_hi (
    .in(Tile_X04_Y0C_hi_unq1),
    .out(Tile_X04_Y0C_hi_out)
);
mantle_wire__typeBit8 Tile_X04_Y0C_lo (
    .in(Tile_X04_Y0C_lo_unq1),
    .out(Tile_X04_Y0C_lo_out)
);
wire [15:0] Tile_X04_Y0C_tile_id_out;
assign Tile_X04_Y0C_tile_id_out = {Tile_X04_Y0C_lo_out[7],Tile_X04_Y0C_lo_out[7:6],Tile_X04_Y0C_lo_out[6:5],Tile_X04_Y0C_hi_out[5],Tile_X04_Y0C_lo_out[4],Tile_X04_Y0C_lo_out[4:3],Tile_X04_Y0C_lo_out[3:2],Tile_X04_Y0C_lo_out[2],Tile_X04_Y0C_hi_out[2:1],Tile_X04_Y0C_lo_out[0],Tile_X04_Y0C_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X04_Y0C_tile_id (
    .in(Tile_X04_Y0C_tile_id_in),
    .out(Tile_X04_Y0C_tile_id_out)
);
Tile_PE Tile_X04_Y0D (
    .SB_T0_EAST_SB_IN_B1(Tile_X05_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X05_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X04_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X04_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X04_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X04_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X04_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X04_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X04_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X04_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X04_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X04_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X03_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X03_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X04_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X04_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X05_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X05_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X04_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X04_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X04_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X04_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X04_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X04_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X04_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X04_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X04_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X04_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X03_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X03_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X04_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X04_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X05_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X05_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X04_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X04_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X04_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X04_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X04_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X04_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X04_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X04_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X04_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X04_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X03_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X03_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X04_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X04_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X05_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X05_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X04_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X04_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X04_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X04_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X04_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X04_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X04_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X04_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X04_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X04_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X03_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X03_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X04_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X04_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X05_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X05_Y0D_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X04_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X04_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X04_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X04_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X04_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X04_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X04_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X04_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X04_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X04_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X03_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X03_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X04_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X04_Y0D_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X04_Y0C_clk_out),
    .clk_out(Tile_X04_Y0D_clk_out),
    .clk_pass_through(Tile_X04_Y0C_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X04_Y0D_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X04_Y0D_clk_pass_through_out_right),
    .config_config_addr(Tile_X04_Y0C_config_out_config_addr),
    .config_config_data(Tile_X04_Y0C_config_out_config_data),
    .config_out_config_addr(Tile_X04_Y0D_config_out_config_addr),
    .config_out_config_data(Tile_X04_Y0D_config_out_config_data),
    .config_out_read(Tile_X04_Y0D_config_out_read),
    .config_out_write(Tile_X04_Y0D_config_out_write),
    .config_read(Tile_X04_Y0C_config_out_read),
    .config_write(Tile_X04_Y0C_config_out_write),
    .hi(Tile_X04_Y0D_hi_unq1),
    .lo(Tile_X04_Y0D_lo_unq1),
    .read_config_data(Tile_X04_Y0D_read_config_data),
    .read_config_data_in(Tile_X04_Y0C_read_config_data),
    .reset(Tile_X04_Y0C_reset_out),
    .reset_out(Tile_X04_Y0D_reset_out),
    .stall(Tile_X04_Y0C_stall_out),
    .stall_out(Tile_X04_Y0D_stall_out),
    .tile_id(Tile_X04_Y0D_tile_id_in)
);
mantle_wire__typeBit9 Tile_X04_Y0D_hi (
    .in(Tile_X04_Y0D_hi_unq1),
    .out(Tile_X04_Y0D_hi_out)
);
mantle_wire__typeBit8 Tile_X04_Y0D_lo (
    .in(Tile_X04_Y0D_lo_unq1),
    .out(Tile_X04_Y0D_lo_out)
);
wire [15:0] Tile_X04_Y0D_tile_id_out;
assign Tile_X04_Y0D_tile_id_out = {Tile_X04_Y0D_lo_out[7],Tile_X04_Y0D_lo_out[7:6],Tile_X04_Y0D_lo_out[6:5],Tile_X04_Y0D_hi_out[5],Tile_X04_Y0D_lo_out[4],Tile_X04_Y0D_lo_out[4:3],Tile_X04_Y0D_lo_out[3:2],Tile_X04_Y0D_lo_out[2],Tile_X04_Y0D_hi_out[2:1],Tile_X04_Y0D_lo_out[0],Tile_X04_Y0D_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X04_Y0D_tile_id (
    .in(Tile_X04_Y0D_tile_id_in),
    .out(Tile_X04_Y0D_tile_id_out)
);
Tile_PE Tile_X04_Y0E (
    .SB_T0_EAST_SB_IN_B1(Tile_X05_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X05_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X04_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X04_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X04_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X04_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X04_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X04_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X04_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X04_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X04_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X04_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X03_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X03_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X04_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X04_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X05_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X05_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X04_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X04_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X04_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X04_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X04_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X04_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X04_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X04_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X04_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X04_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X03_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X03_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X04_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X04_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X05_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X05_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X04_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X04_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X04_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X04_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X04_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X04_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X04_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X04_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X04_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X04_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X03_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X03_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X04_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X04_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X05_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X05_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X04_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X04_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X04_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X04_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X04_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X04_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X04_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X04_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X04_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X04_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X03_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X03_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X04_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X04_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X05_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X05_Y0E_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X04_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X04_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X04_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X04_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X04_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X04_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X04_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X04_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X04_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X04_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X03_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X03_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X04_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X04_Y0E_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X04_Y0D_clk_out),
    .clk_out(Tile_X04_Y0E_clk_out),
    .clk_pass_through(Tile_X04_Y0D_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X04_Y0E_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X04_Y0E_clk_pass_through_out_right),
    .config_config_addr(Tile_X04_Y0D_config_out_config_addr),
    .config_config_data(Tile_X04_Y0D_config_out_config_data),
    .config_out_config_addr(Tile_X04_Y0E_config_out_config_addr),
    .config_out_config_data(Tile_X04_Y0E_config_out_config_data),
    .config_out_read(Tile_X04_Y0E_config_out_read),
    .config_out_write(Tile_X04_Y0E_config_out_write),
    .config_read(Tile_X04_Y0D_config_out_read),
    .config_write(Tile_X04_Y0D_config_out_write),
    .hi(Tile_X04_Y0E_hi_unq1),
    .lo(Tile_X04_Y0E_lo_unq1),
    .read_config_data(Tile_X04_Y0E_read_config_data),
    .read_config_data_in(Tile_X04_Y0D_read_config_data),
    .reset(Tile_X04_Y0D_reset_out),
    .reset_out(Tile_X04_Y0E_reset_out),
    .stall(Tile_X04_Y0D_stall_out),
    .stall_out(Tile_X04_Y0E_stall_out),
    .tile_id(Tile_X04_Y0E_tile_id_in)
);
mantle_wire__typeBit9 Tile_X04_Y0E_hi (
    .in(Tile_X04_Y0E_hi_unq1),
    .out(Tile_X04_Y0E_hi_out)
);
mantle_wire__typeBit8 Tile_X04_Y0E_lo (
    .in(Tile_X04_Y0E_lo_unq1),
    .out(Tile_X04_Y0E_lo_out)
);
wire [15:0] Tile_X04_Y0E_tile_id_out;
assign Tile_X04_Y0E_tile_id_out = {Tile_X04_Y0E_lo_out[7],Tile_X04_Y0E_lo_out[7:6],Tile_X04_Y0E_lo_out[6:5],Tile_X04_Y0E_hi_out[5],Tile_X04_Y0E_lo_out[4],Tile_X04_Y0E_lo_out[4:3],Tile_X04_Y0E_lo_out[3:2],Tile_X04_Y0E_lo_out[2],Tile_X04_Y0E_hi_out[2:1],Tile_X04_Y0E_hi_out[1],Tile_X04_Y0E_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X04_Y0E_tile_id (
    .in(Tile_X04_Y0E_tile_id_in),
    .out(Tile_X04_Y0E_tile_id_out)
);
Tile_PE Tile_X04_Y0F (
    .SB_T0_EAST_SB_IN_B1(Tile_X05_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X05_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X04_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X04_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X04_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X04_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X04_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X04_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X04_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X04_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X04_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X04_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X03_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X03_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X04_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X04_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X05_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X05_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X04_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X04_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X04_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X04_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X04_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X04_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X04_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X04_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X04_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X04_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X03_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X03_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X04_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X04_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X05_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X05_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X04_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X04_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X04_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X04_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X04_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X04_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X04_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X04_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X04_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X04_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X03_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X03_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X04_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X04_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X05_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X05_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X04_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X04_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X04_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X04_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X04_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X04_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X04_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X04_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X04_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X04_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X03_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X03_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X04_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X04_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X05_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X05_Y0F_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X04_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X04_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X04_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X04_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X04_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X04_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X04_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X04_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X04_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X04_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X03_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X03_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X04_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X04_Y0F_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X04_Y0E_clk_out),
    .clk_out(Tile_X04_Y0F_clk_out),
    .clk_pass_through(Tile_X04_Y0E_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X04_Y0F_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X04_Y0F_clk_pass_through_out_right),
    .config_config_addr(Tile_X04_Y0E_config_out_config_addr),
    .config_config_data(Tile_X04_Y0E_config_out_config_data),
    .config_out_config_addr(Tile_X04_Y0F_config_out_config_addr),
    .config_out_config_data(Tile_X04_Y0F_config_out_config_data),
    .config_out_read(Tile_X04_Y0F_config_out_read),
    .config_out_write(Tile_X04_Y0F_config_out_write),
    .config_read(Tile_X04_Y0E_config_out_read),
    .config_write(Tile_X04_Y0E_config_out_write),
    .hi(Tile_X04_Y0F_hi_unq1),
    .lo(Tile_X04_Y0F_lo_unq1),
    .read_config_data(Tile_X04_Y0F_read_config_data),
    .read_config_data_in(Tile_X04_Y0E_read_config_data),
    .reset(Tile_X04_Y0E_reset_out),
    .reset_out(Tile_X04_Y0F_reset_out),
    .stall(Tile_X04_Y0E_stall_out),
    .stall_out(Tile_X04_Y0F_stall_out),
    .tile_id(Tile_X04_Y0F_tile_id_in)
);
mantle_wire__typeBit9 Tile_X04_Y0F_hi (
    .in(Tile_X04_Y0F_hi_unq1),
    .out(Tile_X04_Y0F_hi_out)
);
mantle_wire__typeBit8 Tile_X04_Y0F_lo (
    .in(Tile_X04_Y0F_lo_unq1),
    .out(Tile_X04_Y0F_lo_out)
);
wire [15:0] Tile_X04_Y0F_tile_id_out;
assign Tile_X04_Y0F_tile_id_out = {Tile_X04_Y0F_lo_out[7],Tile_X04_Y0F_lo_out[7:6],Tile_X04_Y0F_lo_out[6:5],Tile_X04_Y0F_hi_out[5],Tile_X04_Y0F_lo_out[4],Tile_X04_Y0F_lo_out[4:3],Tile_X04_Y0F_lo_out[3:2],Tile_X04_Y0F_lo_out[2],Tile_X04_Y0F_hi_out[2:1],Tile_X04_Y0F_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X04_Y0F_tile_id (
    .in(Tile_X04_Y0F_tile_id_in),
    .out(Tile_X04_Y0F_tile_id_out)
);
Tile_PE Tile_X04_Y10 (
    .SB_T0_EAST_SB_IN_B1(Tile_X05_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X05_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X04_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X04_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X04_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X04_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X04_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X04_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T0_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X04_Y10_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X04_Y10_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X03_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X03_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X04_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X04_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X05_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X05_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X04_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X04_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X04_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X04_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X04_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X04_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T1_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X04_Y10_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X04_Y10_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X03_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X03_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X04_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X04_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X05_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X05_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X04_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X04_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X04_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X04_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X04_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X04_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T2_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X04_Y10_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X04_Y10_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X03_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X03_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X04_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X04_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X05_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X05_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X04_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X04_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X04_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X04_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X04_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X04_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T3_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X04_Y10_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X04_Y10_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X03_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X03_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X04_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X04_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X05_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X05_Y10_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X04_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X04_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X04_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X04_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X04_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X04_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T4_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X04_Y10_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X04_Y10_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X03_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X03_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X04_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X04_Y10_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X04_Y0F_clk_out),
    .clk_out(Tile_X04_Y10_clk_out),
    .clk_pass_through(Tile_X04_Y0F_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X04_Y10_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X04_Y10_clk_pass_through_out_right),
    .config_config_addr(Tile_X04_Y0F_config_out_config_addr),
    .config_config_data(Tile_X04_Y0F_config_out_config_data),
    .config_out_config_addr(Tile_X04_Y10_config_out_config_addr),
    .config_out_config_data(Tile_X04_Y10_config_out_config_data),
    .config_out_read(Tile_X04_Y10_config_out_read),
    .config_out_write(Tile_X04_Y10_config_out_write),
    .config_read(Tile_X04_Y0F_config_out_read),
    .config_write(Tile_X04_Y0F_config_out_write),
    .hi(Tile_X04_Y10_hi),
    .lo(Tile_X04_Y10_lo_unq1),
    .read_config_data(Tile_X04_Y10_read_config_data),
    .read_config_data_in(Tile_X04_Y0F_read_config_data),
    .reset(Tile_X04_Y0F_reset_out),
    .reset_out(Tile_X04_Y10_reset_out),
    .stall(Tile_X04_Y0F_stall_out),
    .stall_out(Tile_X04_Y10_stall_out),
    .tile_id(Tile_X04_Y10_tile_id_in)
);
mantle_wire__typeBit8 Tile_X04_Y10_lo (
    .in(Tile_X04_Y10_lo_unq1),
    .out(Tile_X04_Y10_lo_out)
);
wire [15:0] Tile_X04_Y10_tile_id_out;
assign Tile_X04_Y10_tile_id_out = {Tile_X04_Y10_lo_out[7],Tile_X04_Y10_lo_out[7:6],Tile_X04_Y10_lo_out[6:5],Tile_X04_Y10_hi[5],Tile_X04_Y10_lo_out[4],Tile_X04_Y10_lo_out[4:3],Tile_X04_Y10_lo_out[3:2],Tile_X04_Y10_hi[2],Tile_X04_Y10_lo_out[1],Tile_X04_Y10_lo_out[1:0],Tile_X04_Y10_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X04_Y10_tile_id (
    .in(Tile_X04_Y10_tile_id_in),
    .out(Tile_X04_Y10_tile_id_out)
);
wire [15:0] Tile_X05_Y00_tile_id;
assign Tile_X05_Y00_tile_id = {Tile_X05_Y00_lo[7],Tile_X05_Y00_lo[7:6],Tile_X05_Y00_lo[6:5],Tile_X05_Y00_hi[5],Tile_X05_Y00_lo[4],Tile_X05_Y00_hi[4],Tile_X05_Y00_lo[3],Tile_X05_Y00_lo[3:2],Tile_X05_Y00_lo[2:1],Tile_X05_Y00_lo[1:0],Tile_X05_Y00_lo[0]};
Tile_io_core Tile_X05_Y00 (
    .tile_id(Tile_X05_Y00_tile_id),
    .glb2io_1(glb2io_1_X05_Y00),
    .f2io_1(Tile_X05_Y01_SB_T0_NORTH_SB_OUT_B1),
    .io2glb_1(Tile_X05_Y00_io2glb_1),
    .io2f_1(Tile_X05_Y00_io2f_1),
    .glb2io_16(glb2io_16_X05_Y00),
    .f2io_16(Tile_X05_Y01_SB_T0_NORTH_SB_OUT_B16),
    .io2glb_16(Tile_X05_Y00_io2glb_16),
    .io2f_16(Tile_X05_Y00_io2f_16),
    .hi(Tile_X05_Y00_hi),
    .lo(Tile_X05_Y00_lo)
);
Tile_PE Tile_X05_Y01 (
    .SB_T0_EAST_SB_IN_B1(Tile_X06_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X06_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X05_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X05_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X05_Y00_io2f_1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X05_Y00_io2f_16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X05_Y01_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X05_Y01_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X05_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X05_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X05_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X05_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X04_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X04_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X05_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X05_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X06_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X06_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X05_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X05_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X05_Y00_io2f_1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X05_Y00_io2f_16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X05_Y01_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X05_Y01_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X05_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X05_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X05_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X05_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X04_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X04_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X05_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X05_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X06_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X06_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X05_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X05_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X05_Y00_io2f_1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X05_Y00_io2f_16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X05_Y01_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X05_Y01_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X05_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X05_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X05_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X05_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X04_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X04_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X05_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X05_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X06_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X06_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X05_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X05_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X05_Y00_io2f_1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X05_Y00_io2f_16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X05_Y01_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X05_Y01_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X05_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X05_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X05_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X05_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X04_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X04_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X05_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X05_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X06_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X06_Y01_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X05_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X05_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X05_Y00_io2f_1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X05_Y00_io2f_16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X05_Y01_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X05_Y01_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X05_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X05_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X05_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X05_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X04_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X04_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X05_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X05_Y01_SB_T4_WEST_SB_OUT_B16),
    .clk(clk),
    .clk_out(Tile_X05_Y01_clk_out),
    .clk_pass_through(clk),
    .clk_pass_through_out_bot(Tile_X05_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X05_Y01_clk_pass_through_out_right),
    .config_config_addr(config_5_config_addr),
    .config_config_data(config_5_config_data),
    .config_out_config_addr(Tile_X05_Y01_config_out_config_addr),
    .config_out_config_data(Tile_X05_Y01_config_out_config_data),
    .config_out_read(Tile_X05_Y01_config_out_read),
    .config_out_write(Tile_X05_Y01_config_out_write),
    .config_read(config_5_read),
    .config_write(config_5_write),
    .hi(Tile_X05_Y01_hi),
    .lo(Tile_X05_Y01_lo_unq1),
    .read_config_data(Tile_X05_Y01_read_config_data),
    .read_config_data_in(const_0_32_out),
    .reset(reset),
    .reset_out(Tile_X05_Y01_reset_out),
    .stall(stall[5]),
    .stall_out(Tile_X05_Y01_stall_out),
    .tile_id(Tile_X05_Y01_tile_id_in)
);
mantle_wire__typeBit8 Tile_X05_Y01_lo (
    .in(Tile_X05_Y01_lo_unq1),
    .out(Tile_X05_Y01_lo_out)
);
wire [15:0] Tile_X05_Y01_tile_id_out;
assign Tile_X05_Y01_tile_id_out = {Tile_X05_Y01_lo_out[7],Tile_X05_Y01_lo_out[7:6],Tile_X05_Y01_lo_out[6:5],Tile_X05_Y01_hi[5],Tile_X05_Y01_lo_out[4],Tile_X05_Y01_hi[4],Tile_X05_Y01_lo_out[3],Tile_X05_Y01_lo_out[3:2],Tile_X05_Y01_lo_out[2:1],Tile_X05_Y01_lo_out[1:0],Tile_X05_Y01_hi[0]};
mantle_wire__typeBitIn16 Tile_X05_Y01_tile_id (
    .in(Tile_X05_Y01_tile_id_in),
    .out(Tile_X05_Y01_tile_id_out)
);
Tile_PE Tile_X05_Y02 (
    .SB_T0_EAST_SB_IN_B1(Tile_X06_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X06_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X05_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X05_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X05_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X05_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X05_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X05_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X05_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X05_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X05_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X05_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X04_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X04_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X05_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X05_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X06_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X06_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X05_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X05_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X05_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X05_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X05_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X05_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X05_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X05_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X05_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X05_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X04_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X04_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X05_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X05_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X06_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X06_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X05_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X05_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X05_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X05_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X05_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X05_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X05_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X05_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X05_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X05_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X04_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X04_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X05_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X05_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X06_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X06_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X05_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X05_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X05_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X05_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X05_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X05_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X05_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X05_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X05_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X05_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X04_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X04_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X05_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X05_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X06_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X06_Y02_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X05_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X05_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X05_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X05_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X05_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X05_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X05_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X05_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X05_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X05_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X04_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X04_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X05_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X05_Y02_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X05_Y01_clk_out),
    .clk_out(Tile_X05_Y02_clk_out),
    .clk_pass_through(Tile_X05_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X05_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X05_Y02_clk_pass_through_out_right),
    .config_config_addr(Tile_X05_Y01_config_out_config_addr),
    .config_config_data(Tile_X05_Y01_config_out_config_data),
    .config_out_config_addr(Tile_X05_Y02_config_out_config_addr),
    .config_out_config_data(Tile_X05_Y02_config_out_config_data),
    .config_out_read(Tile_X05_Y02_config_out_read),
    .config_out_write(Tile_X05_Y02_config_out_write),
    .config_read(Tile_X05_Y01_config_out_read),
    .config_write(Tile_X05_Y01_config_out_write),
    .hi(Tile_X05_Y02_hi),
    .lo(Tile_X05_Y02_lo_unq1),
    .read_config_data(Tile_X05_Y02_read_config_data),
    .read_config_data_in(Tile_X05_Y01_read_config_data),
    .reset(Tile_X05_Y01_reset_out),
    .reset_out(Tile_X05_Y02_reset_out),
    .stall(Tile_X05_Y01_stall_out),
    .stall_out(Tile_X05_Y02_stall_out),
    .tile_id(Tile_X05_Y02_tile_id_in)
);
mantle_wire__typeBit8 Tile_X05_Y02_lo (
    .in(Tile_X05_Y02_lo_unq1),
    .out(Tile_X05_Y02_lo_out)
);
wire [15:0] Tile_X05_Y02_tile_id_out;
assign Tile_X05_Y02_tile_id_out = {Tile_X05_Y02_lo_out[7],Tile_X05_Y02_lo_out[7:6],Tile_X05_Y02_lo_out[6:5],Tile_X05_Y02_hi[5],Tile_X05_Y02_lo_out[4],Tile_X05_Y02_hi[4],Tile_X05_Y02_lo_out[3],Tile_X05_Y02_lo_out[3:2],Tile_X05_Y02_lo_out[2:1],Tile_X05_Y02_lo_out[1],Tile_X05_Y02_hi[1],Tile_X05_Y02_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X05_Y02_tile_id (
    .in(Tile_X05_Y02_tile_id_in),
    .out(Tile_X05_Y02_tile_id_out)
);
Tile_PE Tile_X05_Y03 (
    .SB_T0_EAST_SB_IN_B1(Tile_X06_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X06_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X05_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X05_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X05_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X05_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X05_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X05_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X05_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X05_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X05_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X05_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X04_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X04_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X05_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X05_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X06_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X06_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X05_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X05_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X05_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X05_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X05_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X05_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X05_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X05_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X05_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X05_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X04_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X04_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X05_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X05_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X06_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X06_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X05_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X05_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X05_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X05_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X05_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X05_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X05_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X05_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X05_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X05_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X04_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X04_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X05_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X05_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X06_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X06_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X05_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X05_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X05_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X05_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X05_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X05_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X05_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X05_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X05_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X05_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X04_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X04_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X05_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X05_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X06_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X06_Y03_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X05_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X05_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X05_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X05_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X05_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X05_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X05_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X05_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X05_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X05_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X04_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X04_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X05_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X05_Y03_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X05_Y02_clk_out),
    .clk_out(Tile_X05_Y03_clk_out),
    .clk_pass_through(Tile_X05_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X05_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X05_Y03_clk_pass_through_out_right),
    .config_config_addr(Tile_X05_Y02_config_out_config_addr),
    .config_config_data(Tile_X05_Y02_config_out_config_data),
    .config_out_config_addr(Tile_X05_Y03_config_out_config_addr),
    .config_out_config_data(Tile_X05_Y03_config_out_config_data),
    .config_out_read(Tile_X05_Y03_config_out_read),
    .config_out_write(Tile_X05_Y03_config_out_write),
    .config_read(Tile_X05_Y02_config_out_read),
    .config_write(Tile_X05_Y02_config_out_write),
    .hi(Tile_X05_Y03_hi_unq1),
    .lo(Tile_X05_Y03_lo_unq1),
    .read_config_data(Tile_X05_Y03_read_config_data),
    .read_config_data_in(Tile_X05_Y02_read_config_data),
    .reset(Tile_X05_Y02_reset_out),
    .reset_out(Tile_X05_Y03_reset_out),
    .stall(Tile_X05_Y02_stall_out),
    .stall_out(Tile_X05_Y03_stall_out),
    .tile_id(Tile_X05_Y03_tile_id_in)
);
mantle_wire__typeBit9 Tile_X05_Y03_hi (
    .in(Tile_X05_Y03_hi_unq1),
    .out(Tile_X05_Y03_hi_out)
);
mantle_wire__typeBit8 Tile_X05_Y03_lo (
    .in(Tile_X05_Y03_lo_unq1),
    .out(Tile_X05_Y03_lo_out)
);
wire [15:0] Tile_X05_Y03_tile_id_out;
assign Tile_X05_Y03_tile_id_out = {Tile_X05_Y03_lo_out[7],Tile_X05_Y03_lo_out[7:6],Tile_X05_Y03_lo_out[6:5],Tile_X05_Y03_hi_out[5],Tile_X05_Y03_lo_out[4],Tile_X05_Y03_hi_out[4],Tile_X05_Y03_lo_out[3],Tile_X05_Y03_lo_out[3:2],Tile_X05_Y03_lo_out[2:1],Tile_X05_Y03_lo_out[1],Tile_X05_Y03_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X05_Y03_tile_id (
    .in(Tile_X05_Y03_tile_id_in),
    .out(Tile_X05_Y03_tile_id_out)
);
Tile_PE Tile_X05_Y04 (
    .SB_T0_EAST_SB_IN_B1(Tile_X06_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X06_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X05_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X05_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X05_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X05_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X05_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X05_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X05_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X05_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X05_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X05_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X04_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X04_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X05_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X05_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X06_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X06_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X05_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X05_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X05_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X05_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X05_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X05_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X05_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X05_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X05_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X05_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X04_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X04_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X05_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X05_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X06_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X06_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X05_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X05_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X05_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X05_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X05_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X05_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X05_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X05_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X05_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X05_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X04_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X04_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X05_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X05_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X06_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X06_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X05_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X05_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X05_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X05_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X05_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X05_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X05_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X05_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X05_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X05_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X04_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X04_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X05_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X05_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X06_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X06_Y04_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X05_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X05_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X05_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X05_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X05_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X05_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X05_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X05_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X05_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X05_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X04_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X04_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X05_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X05_Y04_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X05_Y03_clk_out),
    .clk_out(Tile_X05_Y04_clk_out),
    .clk_pass_through(Tile_X05_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X05_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X05_Y04_clk_pass_through_out_right),
    .config_config_addr(Tile_X05_Y03_config_out_config_addr),
    .config_config_data(Tile_X05_Y03_config_out_config_data),
    .config_out_config_addr(Tile_X05_Y04_config_out_config_addr),
    .config_out_config_data(Tile_X05_Y04_config_out_config_data),
    .config_out_read(Tile_X05_Y04_config_out_read),
    .config_out_write(Tile_X05_Y04_config_out_write),
    .config_read(Tile_X05_Y03_config_out_read),
    .config_write(Tile_X05_Y03_config_out_write),
    .hi(Tile_X05_Y04_hi),
    .lo(Tile_X05_Y04_lo_unq1),
    .read_config_data(Tile_X05_Y04_read_config_data),
    .read_config_data_in(Tile_X05_Y03_read_config_data),
    .reset(Tile_X05_Y03_reset_out),
    .reset_out(Tile_X05_Y04_reset_out),
    .stall(Tile_X05_Y03_stall_out),
    .stall_out(Tile_X05_Y04_stall_out),
    .tile_id(Tile_X05_Y04_tile_id_in)
);
mantle_wire__typeBit8 Tile_X05_Y04_lo (
    .in(Tile_X05_Y04_lo_unq1),
    .out(Tile_X05_Y04_lo_out)
);
wire [15:0] Tile_X05_Y04_tile_id_out;
assign Tile_X05_Y04_tile_id_out = {Tile_X05_Y04_lo_out[7],Tile_X05_Y04_lo_out[7:6],Tile_X05_Y04_lo_out[6:5],Tile_X05_Y04_hi[5],Tile_X05_Y04_lo_out[4],Tile_X05_Y04_hi[4],Tile_X05_Y04_lo_out[3],Tile_X05_Y04_lo_out[3:2],Tile_X05_Y04_lo_out[2:1],Tile_X05_Y04_hi[1],Tile_X05_Y04_lo_out[0],Tile_X05_Y04_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X05_Y04_tile_id (
    .in(Tile_X05_Y04_tile_id_in),
    .out(Tile_X05_Y04_tile_id_out)
);
Tile_PE Tile_X05_Y05 (
    .SB_T0_EAST_SB_IN_B1(Tile_X06_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X06_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X05_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X05_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X05_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X05_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X05_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X05_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X05_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X05_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X05_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X05_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X04_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X04_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X05_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X05_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X06_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X06_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X05_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X05_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X05_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X05_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X05_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X05_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X05_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X05_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X05_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X05_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X04_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X04_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X05_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X05_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X06_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X06_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X05_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X05_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X05_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X05_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X05_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X05_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X05_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X05_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X05_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X05_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X04_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X04_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X05_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X05_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X06_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X06_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X05_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X05_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X05_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X05_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X05_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X05_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X05_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X05_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X05_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X05_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X04_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X04_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X05_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X05_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X06_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X06_Y05_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X05_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X05_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X05_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X05_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X05_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X05_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X05_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X05_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X05_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X05_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X04_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X04_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X05_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X05_Y05_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X05_Y04_clk_out),
    .clk_out(Tile_X05_Y05_clk_out),
    .clk_pass_through(Tile_X05_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X05_Y05_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X05_Y05_clk_pass_through_out_right),
    .config_config_addr(Tile_X05_Y04_config_out_config_addr),
    .config_config_data(Tile_X05_Y04_config_out_config_data),
    .config_out_config_addr(Tile_X05_Y05_config_out_config_addr),
    .config_out_config_data(Tile_X05_Y05_config_out_config_data),
    .config_out_read(Tile_X05_Y05_config_out_read),
    .config_out_write(Tile_X05_Y05_config_out_write),
    .config_read(Tile_X05_Y04_config_out_read),
    .config_write(Tile_X05_Y04_config_out_write),
    .hi(Tile_X05_Y05_hi),
    .lo(Tile_X05_Y05_lo_unq1),
    .read_config_data(Tile_X05_Y05_read_config_data),
    .read_config_data_in(Tile_X05_Y04_read_config_data),
    .reset(Tile_X05_Y04_reset_out),
    .reset_out(Tile_X05_Y05_reset_out),
    .stall(Tile_X05_Y04_stall_out),
    .stall_out(Tile_X05_Y05_stall_out),
    .tile_id(Tile_X05_Y05_tile_id_in)
);
mantle_wire__typeBit8 Tile_X05_Y05_lo (
    .in(Tile_X05_Y05_lo_unq1),
    .out(Tile_X05_Y05_lo_out)
);
wire [15:0] Tile_X05_Y05_tile_id_out;
assign Tile_X05_Y05_tile_id_out = {Tile_X05_Y05_lo_out[7],Tile_X05_Y05_lo_out[7:6],Tile_X05_Y05_lo_out[6:5],Tile_X05_Y05_hi[5],Tile_X05_Y05_lo_out[4],Tile_X05_Y05_hi[4],Tile_X05_Y05_lo_out[3],Tile_X05_Y05_lo_out[3:2],Tile_X05_Y05_lo_out[2:1],Tile_X05_Y05_hi[1],Tile_X05_Y05_lo_out[0],Tile_X05_Y05_hi[0]};
mantle_wire__typeBitIn16 Tile_X05_Y05_tile_id (
    .in(Tile_X05_Y05_tile_id_in),
    .out(Tile_X05_Y05_tile_id_out)
);
Tile_PE Tile_X05_Y06 (
    .SB_T0_EAST_SB_IN_B1(Tile_X06_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X06_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X05_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X05_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X05_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X05_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X05_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X05_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X05_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X05_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X05_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X05_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X04_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X04_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X05_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X05_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X06_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X06_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X05_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X05_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X05_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X05_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X05_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X05_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X05_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X05_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X05_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X05_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X04_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X04_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X05_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X05_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X06_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X06_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X05_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X05_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X05_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X05_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X05_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X05_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X05_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X05_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X05_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X05_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X04_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X04_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X05_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X05_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X06_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X06_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X05_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X05_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X05_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X05_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X05_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X05_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X05_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X05_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X05_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X05_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X04_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X04_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X05_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X05_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X06_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X06_Y06_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X05_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X05_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X05_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X05_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X05_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X05_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X05_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X05_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X05_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X05_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X04_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X04_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X05_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X05_Y06_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X05_Y05_clk_out),
    .clk_out(Tile_X05_Y06_clk_out),
    .clk_pass_through(Tile_X05_Y05_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X05_Y06_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X05_Y06_clk_pass_through_out_right),
    .config_config_addr(Tile_X05_Y05_config_out_config_addr),
    .config_config_data(Tile_X05_Y05_config_out_config_data),
    .config_out_config_addr(Tile_X05_Y06_config_out_config_addr),
    .config_out_config_data(Tile_X05_Y06_config_out_config_data),
    .config_out_read(Tile_X05_Y06_config_out_read),
    .config_out_write(Tile_X05_Y06_config_out_write),
    .config_read(Tile_X05_Y05_config_out_read),
    .config_write(Tile_X05_Y05_config_out_write),
    .hi(Tile_X05_Y06_hi),
    .lo(Tile_X05_Y06_lo_unq1),
    .read_config_data(Tile_X05_Y06_read_config_data),
    .read_config_data_in(Tile_X05_Y05_read_config_data),
    .reset(Tile_X05_Y05_reset_out),
    .reset_out(Tile_X05_Y06_reset_out),
    .stall(Tile_X05_Y05_stall_out),
    .stall_out(Tile_X05_Y06_stall_out),
    .tile_id(Tile_X05_Y06_tile_id_in)
);
mantle_wire__typeBit8 Tile_X05_Y06_lo (
    .in(Tile_X05_Y06_lo_unq1),
    .out(Tile_X05_Y06_lo_out)
);
wire [15:0] Tile_X05_Y06_tile_id_out;
assign Tile_X05_Y06_tile_id_out = {Tile_X05_Y06_lo_out[7],Tile_X05_Y06_lo_out[7:6],Tile_X05_Y06_lo_out[6:5],Tile_X05_Y06_hi[5],Tile_X05_Y06_lo_out[4],Tile_X05_Y06_hi[4],Tile_X05_Y06_lo_out[3],Tile_X05_Y06_lo_out[3:2],Tile_X05_Y06_lo_out[2:1],Tile_X05_Y06_hi[1],Tile_X05_Y06_hi[1],Tile_X05_Y06_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X05_Y06_tile_id (
    .in(Tile_X05_Y06_tile_id_in),
    .out(Tile_X05_Y06_tile_id_out)
);
Tile_PE Tile_X05_Y07 (
    .SB_T0_EAST_SB_IN_B1(Tile_X06_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X06_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X05_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X05_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X05_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X05_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X05_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X05_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X05_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X05_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X05_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X05_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X04_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X04_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X05_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X05_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X06_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X06_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X05_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X05_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X05_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X05_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X05_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X05_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X05_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X05_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X05_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X05_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X04_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X04_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X05_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X05_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X06_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X06_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X05_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X05_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X05_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X05_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X05_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X05_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X05_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X05_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X05_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X05_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X04_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X04_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X05_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X05_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X06_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X06_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X05_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X05_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X05_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X05_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X05_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X05_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X05_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X05_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X05_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X05_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X04_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X04_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X05_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X05_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X06_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X06_Y07_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X05_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X05_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X05_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X05_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X05_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X05_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X05_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X05_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X05_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X05_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X04_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X04_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X05_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X05_Y07_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X05_Y06_clk_out),
    .clk_out(Tile_X05_Y07_clk_out),
    .clk_pass_through(Tile_X05_Y06_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X05_Y07_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X05_Y07_clk_pass_through_out_right),
    .config_config_addr(Tile_X05_Y06_config_out_config_addr),
    .config_config_data(Tile_X05_Y06_config_out_config_data),
    .config_out_config_addr(Tile_X05_Y07_config_out_config_addr),
    .config_out_config_data(Tile_X05_Y07_config_out_config_data),
    .config_out_read(Tile_X05_Y07_config_out_read),
    .config_out_write(Tile_X05_Y07_config_out_write),
    .config_read(Tile_X05_Y06_config_out_read),
    .config_write(Tile_X05_Y06_config_out_write),
    .hi(Tile_X05_Y07_hi_unq1),
    .lo(Tile_X05_Y07_lo_unq1),
    .read_config_data(Tile_X05_Y07_read_config_data),
    .read_config_data_in(Tile_X05_Y06_read_config_data),
    .reset(Tile_X05_Y06_reset_out),
    .reset_out(Tile_X05_Y07_reset_out),
    .stall(Tile_X05_Y06_stall_out),
    .stall_out(Tile_X05_Y07_stall_out),
    .tile_id(Tile_X05_Y07_tile_id_in)
);
mantle_wire__typeBit9 Tile_X05_Y07_hi (
    .in(Tile_X05_Y07_hi_unq1),
    .out(Tile_X05_Y07_hi_out)
);
mantle_wire__typeBit8 Tile_X05_Y07_lo (
    .in(Tile_X05_Y07_lo_unq1),
    .out(Tile_X05_Y07_lo_out)
);
wire [15:0] Tile_X05_Y07_tile_id_out;
assign Tile_X05_Y07_tile_id_out = {Tile_X05_Y07_lo_out[7],Tile_X05_Y07_lo_out[7:6],Tile_X05_Y07_lo_out[6:5],Tile_X05_Y07_hi_out[5],Tile_X05_Y07_lo_out[4],Tile_X05_Y07_hi_out[4],Tile_X05_Y07_lo_out[3],Tile_X05_Y07_lo_out[3:2],Tile_X05_Y07_lo_out[2:1],Tile_X05_Y07_hi_out[1],Tile_X05_Y07_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X05_Y07_tile_id (
    .in(Tile_X05_Y07_tile_id_in),
    .out(Tile_X05_Y07_tile_id_out)
);
Tile_PE Tile_X05_Y08 (
    .SB_T0_EAST_SB_IN_B1(Tile_X06_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X06_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X05_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X05_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X05_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X05_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X05_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X05_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X05_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X05_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X05_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X05_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X04_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X04_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X05_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X05_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X06_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X06_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X05_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X05_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X05_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X05_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X05_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X05_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X05_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X05_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X05_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X05_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X04_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X04_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X05_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X05_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X06_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X06_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X05_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X05_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X05_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X05_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X05_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X05_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X05_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X05_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X05_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X05_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X04_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X04_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X05_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X05_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X06_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X06_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X05_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X05_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X05_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X05_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X05_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X05_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X05_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X05_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X05_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X05_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X04_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X04_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X05_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X05_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X06_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X06_Y08_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X05_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X05_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X05_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X05_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X05_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X05_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X05_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X05_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X05_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X05_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X04_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X04_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X05_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X05_Y08_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X05_Y07_clk_out),
    .clk_out(Tile_X05_Y08_clk_out),
    .clk_pass_through(Tile_X05_Y07_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X05_Y08_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X05_Y08_clk_pass_through_out_right),
    .config_config_addr(Tile_X05_Y07_config_out_config_addr),
    .config_config_data(Tile_X05_Y07_config_out_config_data),
    .config_out_config_addr(Tile_X05_Y08_config_out_config_addr),
    .config_out_config_data(Tile_X05_Y08_config_out_config_data),
    .config_out_read(Tile_X05_Y08_config_out_read),
    .config_out_write(Tile_X05_Y08_config_out_write),
    .config_read(Tile_X05_Y07_config_out_read),
    .config_write(Tile_X05_Y07_config_out_write),
    .hi(Tile_X05_Y08_hi),
    .lo(Tile_X05_Y08_lo_unq1),
    .read_config_data(Tile_X05_Y08_read_config_data),
    .read_config_data_in(Tile_X05_Y07_read_config_data),
    .reset(Tile_X05_Y07_reset_out),
    .reset_out(Tile_X05_Y08_reset_out),
    .stall(Tile_X05_Y07_stall_out),
    .stall_out(Tile_X05_Y08_stall_out),
    .tile_id(Tile_X05_Y08_tile_id_in)
);
mantle_wire__typeBit8 Tile_X05_Y08_lo (
    .in(Tile_X05_Y08_lo_unq1),
    .out(Tile_X05_Y08_lo_out)
);
wire [15:0] Tile_X05_Y08_tile_id_out;
assign Tile_X05_Y08_tile_id_out = {Tile_X05_Y08_lo_out[7],Tile_X05_Y08_lo_out[7:6],Tile_X05_Y08_lo_out[6:5],Tile_X05_Y08_hi[5],Tile_X05_Y08_lo_out[4],Tile_X05_Y08_hi[4],Tile_X05_Y08_lo_out[3],Tile_X05_Y08_lo_out[3:2],Tile_X05_Y08_lo_out[2],Tile_X05_Y08_hi[2],Tile_X05_Y08_lo_out[1:0],Tile_X05_Y08_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X05_Y08_tile_id (
    .in(Tile_X05_Y08_tile_id_in),
    .out(Tile_X05_Y08_tile_id_out)
);
Tile_PE Tile_X05_Y09 (
    .SB_T0_EAST_SB_IN_B1(Tile_X06_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X06_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X05_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X05_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X05_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X05_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X05_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X05_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X05_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X05_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X05_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X05_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X04_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X04_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X05_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X05_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X06_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X06_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X05_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X05_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X05_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X05_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X05_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X05_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X05_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X05_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X05_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X05_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X04_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X04_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X05_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X05_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X06_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X06_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X05_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X05_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X05_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X05_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X05_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X05_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X05_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X05_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X05_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X05_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X04_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X04_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X05_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X05_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X06_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X06_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X05_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X05_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X05_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X05_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X05_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X05_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X05_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X05_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X05_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X05_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X04_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X04_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X05_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X05_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X06_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X06_Y09_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X05_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X05_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X05_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X05_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X05_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X05_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X05_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X05_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X05_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X05_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X04_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X04_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X05_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X05_Y09_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X05_Y08_clk_out),
    .clk_out(Tile_X05_Y09_clk_out),
    .clk_pass_through(Tile_X05_Y08_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X05_Y09_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X05_Y09_clk_pass_through_out_right),
    .config_config_addr(ConfigPipeStage_inst5_config_out_config_addr),
    .config_config_data(ConfigPipeStage_inst5_config_out_config_data),
    .config_out_config_addr(Tile_X05_Y09_config_out_config_addr),
    .config_out_config_data(Tile_X05_Y09_config_out_config_data),
    .config_out_read(Tile_X05_Y09_config_out_read),
    .config_out_write(Tile_X05_Y09_config_out_write),
    .config_read(ConfigPipeStage_inst5_config_out_read),
    .config_write(ConfigPipeStage_inst5_config_out_write),
    .hi(Tile_X05_Y09_hi),
    .lo(Tile_X05_Y09_lo_unq1),
    .read_config_data(Tile_X05_Y09_read_config_data),
    .read_config_data_in(Tile_X05_Y08_read_config_data),
    .reset(Tile_X05_Y08_reset_out),
    .reset_out(Tile_X05_Y09_reset_out),
    .stall(Tile_X05_Y08_stall_out),
    .stall_out(Tile_X05_Y09_stall_out),
    .tile_id(Tile_X05_Y09_tile_id_in)
);
mantle_wire__typeBit8 Tile_X05_Y09_lo (
    .in(Tile_X05_Y09_lo_unq1),
    .out(Tile_X05_Y09_lo_out)
);
wire [15:0] Tile_X05_Y09_tile_id_out;
assign Tile_X05_Y09_tile_id_out = {Tile_X05_Y09_lo_out[7],Tile_X05_Y09_lo_out[7:6],Tile_X05_Y09_lo_out[6:5],Tile_X05_Y09_hi[5],Tile_X05_Y09_lo_out[4],Tile_X05_Y09_hi[4],Tile_X05_Y09_lo_out[3],Tile_X05_Y09_lo_out[3:2],Tile_X05_Y09_lo_out[2],Tile_X05_Y09_hi[2],Tile_X05_Y09_lo_out[1:0],Tile_X05_Y09_hi[0]};
mantle_wire__typeBitIn16 Tile_X05_Y09_tile_id (
    .in(Tile_X05_Y09_tile_id_in),
    .out(Tile_X05_Y09_tile_id_out)
);
Tile_PE Tile_X05_Y0A (
    .SB_T0_EAST_SB_IN_B1(Tile_X06_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X06_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X05_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X05_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X05_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X05_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X05_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X05_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X05_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X05_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X05_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X05_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X04_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X04_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X05_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X05_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X06_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X06_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X05_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X05_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X05_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X05_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X05_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X05_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X05_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X05_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X05_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X05_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X04_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X04_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X05_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X05_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X06_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X06_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X05_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X05_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X05_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X05_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X05_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X05_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X05_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X05_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X05_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X05_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X04_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X04_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X05_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X05_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X06_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X06_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X05_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X05_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X05_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X05_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X05_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X05_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X05_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X05_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X05_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X05_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X04_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X04_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X05_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X05_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X06_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X06_Y0A_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X05_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X05_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X05_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X05_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X05_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X05_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X05_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X05_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X05_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X05_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X04_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X04_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X05_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X05_Y0A_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X05_Y09_clk_out),
    .clk_out(Tile_X05_Y0A_clk_out),
    .clk_pass_through(Tile_X05_Y09_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X05_Y0A_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X05_Y0A_clk_pass_through_out_right),
    .config_config_addr(Tile_X05_Y09_config_out_config_addr),
    .config_config_data(Tile_X05_Y09_config_out_config_data),
    .config_out_config_addr(Tile_X05_Y0A_config_out_config_addr),
    .config_out_config_data(Tile_X05_Y0A_config_out_config_data),
    .config_out_read(Tile_X05_Y0A_config_out_read),
    .config_out_write(Tile_X05_Y0A_config_out_write),
    .config_read(Tile_X05_Y09_config_out_read),
    .config_write(Tile_X05_Y09_config_out_write),
    .hi(Tile_X05_Y0A_hi),
    .lo(Tile_X05_Y0A_lo_unq1),
    .read_config_data(Tile_X05_Y0A_read_config_data),
    .read_config_data_in(Tile_X05_Y09_read_config_data),
    .reset(Tile_X05_Y09_reset_out),
    .reset_out(Tile_X05_Y0A_reset_out),
    .stall(Tile_X05_Y09_stall_out),
    .stall_out(Tile_X05_Y0A_stall_out),
    .tile_id(Tile_X05_Y0A_tile_id_in)
);
mantle_wire__typeBit8 Tile_X05_Y0A_lo (
    .in(Tile_X05_Y0A_lo_unq1),
    .out(Tile_X05_Y0A_lo_out)
);
wire [15:0] Tile_X05_Y0A_tile_id_out;
assign Tile_X05_Y0A_tile_id_out = {Tile_X05_Y0A_lo_out[7],Tile_X05_Y0A_lo_out[7:6],Tile_X05_Y0A_lo_out[6:5],Tile_X05_Y0A_hi[5],Tile_X05_Y0A_lo_out[4],Tile_X05_Y0A_hi[4],Tile_X05_Y0A_lo_out[3],Tile_X05_Y0A_lo_out[3:2],Tile_X05_Y0A_lo_out[2],Tile_X05_Y0A_hi[2],Tile_X05_Y0A_lo_out[1],Tile_X05_Y0A_hi[1],Tile_X05_Y0A_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X05_Y0A_tile_id (
    .in(Tile_X05_Y0A_tile_id_in),
    .out(Tile_X05_Y0A_tile_id_out)
);
Tile_PE Tile_X05_Y0B (
    .SB_T0_EAST_SB_IN_B1(Tile_X06_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X06_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X05_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X05_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X05_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X05_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X05_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X05_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X05_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X05_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X05_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X05_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X04_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X04_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X05_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X05_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X06_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X06_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X05_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X05_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X05_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X05_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X05_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X05_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X05_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X05_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X05_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X05_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X04_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X04_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X05_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X05_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X06_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X06_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X05_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X05_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X05_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X05_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X05_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X05_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X05_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X05_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X05_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X05_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X04_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X04_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X05_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X05_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X06_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X06_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X05_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X05_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X05_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X05_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X05_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X05_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X05_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X05_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X05_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X05_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X04_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X04_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X05_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X05_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X06_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X06_Y0B_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X05_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X05_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X05_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X05_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X05_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X05_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X05_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X05_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X05_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X05_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X04_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X04_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X05_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X05_Y0B_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X05_Y0A_clk_out),
    .clk_out(Tile_X05_Y0B_clk_out),
    .clk_pass_through(Tile_X05_Y0A_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X05_Y0B_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X05_Y0B_clk_pass_through_out_right),
    .config_config_addr(Tile_X05_Y0A_config_out_config_addr),
    .config_config_data(Tile_X05_Y0A_config_out_config_data),
    .config_out_config_addr(Tile_X05_Y0B_config_out_config_addr),
    .config_out_config_data(Tile_X05_Y0B_config_out_config_data),
    .config_out_read(Tile_X05_Y0B_config_out_read),
    .config_out_write(Tile_X05_Y0B_config_out_write),
    .config_read(Tile_X05_Y0A_config_out_read),
    .config_write(Tile_X05_Y0A_config_out_write),
    .hi(Tile_X05_Y0B_hi_unq1),
    .lo(Tile_X05_Y0B_lo_unq1),
    .read_config_data(Tile_X05_Y0B_read_config_data),
    .read_config_data_in(Tile_X05_Y0A_read_config_data),
    .reset(Tile_X05_Y0A_reset_out),
    .reset_out(Tile_X05_Y0B_reset_out),
    .stall(Tile_X05_Y0A_stall_out),
    .stall_out(Tile_X05_Y0B_stall_out),
    .tile_id(Tile_X05_Y0B_tile_id_in)
);
mantle_wire__typeBit9 Tile_X05_Y0B_hi (
    .in(Tile_X05_Y0B_hi_unq1),
    .out(Tile_X05_Y0B_hi_out)
);
mantle_wire__typeBit8 Tile_X05_Y0B_lo (
    .in(Tile_X05_Y0B_lo_unq1),
    .out(Tile_X05_Y0B_lo_out)
);
wire [15:0] Tile_X05_Y0B_tile_id_out;
assign Tile_X05_Y0B_tile_id_out = {Tile_X05_Y0B_lo_out[7],Tile_X05_Y0B_lo_out[7:6],Tile_X05_Y0B_lo_out[6:5],Tile_X05_Y0B_hi_out[5],Tile_X05_Y0B_lo_out[4],Tile_X05_Y0B_hi_out[4],Tile_X05_Y0B_lo_out[3],Tile_X05_Y0B_lo_out[3:2],Tile_X05_Y0B_lo_out[2],Tile_X05_Y0B_hi_out[2],Tile_X05_Y0B_lo_out[1],Tile_X05_Y0B_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X05_Y0B_tile_id (
    .in(Tile_X05_Y0B_tile_id_in),
    .out(Tile_X05_Y0B_tile_id_out)
);
Tile_PE Tile_X05_Y0C (
    .SB_T0_EAST_SB_IN_B1(Tile_X06_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X06_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X05_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X05_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X05_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X05_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X05_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X05_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X05_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X05_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X05_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X05_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X04_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X04_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X05_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X05_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X06_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X06_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X05_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X05_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X05_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X05_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X05_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X05_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X05_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X05_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X05_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X05_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X04_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X04_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X05_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X05_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X06_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X06_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X05_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X05_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X05_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X05_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X05_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X05_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X05_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X05_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X05_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X05_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X04_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X04_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X05_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X05_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X06_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X06_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X05_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X05_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X05_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X05_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X05_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X05_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X05_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X05_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X05_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X05_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X04_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X04_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X05_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X05_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X06_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X06_Y0C_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X05_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X05_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X05_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X05_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X05_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X05_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X05_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X05_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X05_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X05_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X04_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X04_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X05_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X05_Y0C_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X05_Y0B_clk_out),
    .clk_out(Tile_X05_Y0C_clk_out),
    .clk_pass_through(Tile_X05_Y0B_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X05_Y0C_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X05_Y0C_clk_pass_through_out_right),
    .config_config_addr(Tile_X05_Y0B_config_out_config_addr),
    .config_config_data(Tile_X05_Y0B_config_out_config_data),
    .config_out_config_addr(Tile_X05_Y0C_config_out_config_addr),
    .config_out_config_data(Tile_X05_Y0C_config_out_config_data),
    .config_out_read(Tile_X05_Y0C_config_out_read),
    .config_out_write(Tile_X05_Y0C_config_out_write),
    .config_read(Tile_X05_Y0B_config_out_read),
    .config_write(Tile_X05_Y0B_config_out_write),
    .hi(Tile_X05_Y0C_hi_unq1),
    .lo(Tile_X05_Y0C_lo_unq1),
    .read_config_data(Tile_X05_Y0C_read_config_data),
    .read_config_data_in(Tile_X05_Y0B_read_config_data),
    .reset(Tile_X05_Y0B_reset_out),
    .reset_out(Tile_X05_Y0C_reset_out),
    .stall(Tile_X05_Y0B_stall_out),
    .stall_out(Tile_X05_Y0C_stall_out),
    .tile_id(Tile_X05_Y0C_tile_id_in)
);
mantle_wire__typeBit9 Tile_X05_Y0C_hi (
    .in(Tile_X05_Y0C_hi_unq1),
    .out(Tile_X05_Y0C_hi_out)
);
mantle_wire__typeBit8 Tile_X05_Y0C_lo (
    .in(Tile_X05_Y0C_lo_unq1),
    .out(Tile_X05_Y0C_lo_out)
);
wire [15:0] Tile_X05_Y0C_tile_id_out;
assign Tile_X05_Y0C_tile_id_out = {Tile_X05_Y0C_lo_out[7],Tile_X05_Y0C_lo_out[7:6],Tile_X05_Y0C_lo_out[6:5],Tile_X05_Y0C_hi_out[5],Tile_X05_Y0C_lo_out[4],Tile_X05_Y0C_hi_out[4],Tile_X05_Y0C_lo_out[3],Tile_X05_Y0C_lo_out[3:2],Tile_X05_Y0C_lo_out[2],Tile_X05_Y0C_hi_out[2:1],Tile_X05_Y0C_lo_out[0],Tile_X05_Y0C_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X05_Y0C_tile_id (
    .in(Tile_X05_Y0C_tile_id_in),
    .out(Tile_X05_Y0C_tile_id_out)
);
Tile_PE Tile_X05_Y0D (
    .SB_T0_EAST_SB_IN_B1(Tile_X06_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X06_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X05_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X05_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X05_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X05_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X05_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X05_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X05_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X05_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X05_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X05_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X04_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X04_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X05_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X05_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X06_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X06_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X05_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X05_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X05_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X05_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X05_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X05_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X05_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X05_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X05_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X05_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X04_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X04_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X05_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X05_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X06_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X06_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X05_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X05_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X05_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X05_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X05_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X05_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X05_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X05_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X05_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X05_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X04_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X04_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X05_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X05_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X06_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X06_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X05_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X05_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X05_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X05_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X05_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X05_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X05_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X05_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X05_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X05_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X04_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X04_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X05_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X05_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X06_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X06_Y0D_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X05_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X05_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X05_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X05_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X05_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X05_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X05_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X05_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X05_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X05_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X04_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X04_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X05_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X05_Y0D_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X05_Y0C_clk_out),
    .clk_out(Tile_X05_Y0D_clk_out),
    .clk_pass_through(Tile_X05_Y0C_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X05_Y0D_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X05_Y0D_clk_pass_through_out_right),
    .config_config_addr(Tile_X05_Y0C_config_out_config_addr),
    .config_config_data(Tile_X05_Y0C_config_out_config_data),
    .config_out_config_addr(Tile_X05_Y0D_config_out_config_addr),
    .config_out_config_data(Tile_X05_Y0D_config_out_config_data),
    .config_out_read(Tile_X05_Y0D_config_out_read),
    .config_out_write(Tile_X05_Y0D_config_out_write),
    .config_read(Tile_X05_Y0C_config_out_read),
    .config_write(Tile_X05_Y0C_config_out_write),
    .hi(Tile_X05_Y0D_hi_unq1),
    .lo(Tile_X05_Y0D_lo_unq1),
    .read_config_data(Tile_X05_Y0D_read_config_data),
    .read_config_data_in(Tile_X05_Y0C_read_config_data),
    .reset(Tile_X05_Y0C_reset_out),
    .reset_out(Tile_X05_Y0D_reset_out),
    .stall(Tile_X05_Y0C_stall_out),
    .stall_out(Tile_X05_Y0D_stall_out),
    .tile_id(Tile_X05_Y0D_tile_id_in)
);
mantle_wire__typeBit9 Tile_X05_Y0D_hi (
    .in(Tile_X05_Y0D_hi_unq1),
    .out(Tile_X05_Y0D_hi_out)
);
mantle_wire__typeBit8 Tile_X05_Y0D_lo (
    .in(Tile_X05_Y0D_lo_unq1),
    .out(Tile_X05_Y0D_lo_out)
);
wire [15:0] Tile_X05_Y0D_tile_id_out;
assign Tile_X05_Y0D_tile_id_out = {Tile_X05_Y0D_lo_out[7],Tile_X05_Y0D_lo_out[7:6],Tile_X05_Y0D_lo_out[6:5],Tile_X05_Y0D_hi_out[5],Tile_X05_Y0D_lo_out[4],Tile_X05_Y0D_hi_out[4],Tile_X05_Y0D_lo_out[3],Tile_X05_Y0D_lo_out[3:2],Tile_X05_Y0D_lo_out[2],Tile_X05_Y0D_hi_out[2:1],Tile_X05_Y0D_lo_out[0],Tile_X05_Y0D_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X05_Y0D_tile_id (
    .in(Tile_X05_Y0D_tile_id_in),
    .out(Tile_X05_Y0D_tile_id_out)
);
Tile_PE Tile_X05_Y0E (
    .SB_T0_EAST_SB_IN_B1(Tile_X06_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X06_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X05_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X05_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X05_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X05_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X05_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X05_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X05_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X05_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X05_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X05_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X04_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X04_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X05_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X05_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X06_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X06_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X05_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X05_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X05_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X05_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X05_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X05_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X05_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X05_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X05_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X05_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X04_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X04_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X05_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X05_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X06_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X06_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X05_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X05_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X05_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X05_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X05_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X05_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X05_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X05_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X05_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X05_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X04_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X04_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X05_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X05_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X06_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X06_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X05_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X05_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X05_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X05_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X05_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X05_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X05_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X05_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X05_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X05_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X04_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X04_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X05_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X05_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X06_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X06_Y0E_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X05_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X05_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X05_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X05_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X05_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X05_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X05_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X05_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X05_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X05_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X04_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X04_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X05_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X05_Y0E_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X05_Y0D_clk_out),
    .clk_out(Tile_X05_Y0E_clk_out),
    .clk_pass_through(Tile_X05_Y0D_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X05_Y0E_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X05_Y0E_clk_pass_through_out_right),
    .config_config_addr(Tile_X05_Y0D_config_out_config_addr),
    .config_config_data(Tile_X05_Y0D_config_out_config_data),
    .config_out_config_addr(Tile_X05_Y0E_config_out_config_addr),
    .config_out_config_data(Tile_X05_Y0E_config_out_config_data),
    .config_out_read(Tile_X05_Y0E_config_out_read),
    .config_out_write(Tile_X05_Y0E_config_out_write),
    .config_read(Tile_X05_Y0D_config_out_read),
    .config_write(Tile_X05_Y0D_config_out_write),
    .hi(Tile_X05_Y0E_hi_unq1),
    .lo(Tile_X05_Y0E_lo_unq1),
    .read_config_data(Tile_X05_Y0E_read_config_data),
    .read_config_data_in(Tile_X05_Y0D_read_config_data),
    .reset(Tile_X05_Y0D_reset_out),
    .reset_out(Tile_X05_Y0E_reset_out),
    .stall(Tile_X05_Y0D_stall_out),
    .stall_out(Tile_X05_Y0E_stall_out),
    .tile_id(Tile_X05_Y0E_tile_id_in)
);
mantle_wire__typeBit9 Tile_X05_Y0E_hi (
    .in(Tile_X05_Y0E_hi_unq1),
    .out(Tile_X05_Y0E_hi_out)
);
mantle_wire__typeBit8 Tile_X05_Y0E_lo (
    .in(Tile_X05_Y0E_lo_unq1),
    .out(Tile_X05_Y0E_lo_out)
);
wire [15:0] Tile_X05_Y0E_tile_id_out;
assign Tile_X05_Y0E_tile_id_out = {Tile_X05_Y0E_lo_out[7],Tile_X05_Y0E_lo_out[7:6],Tile_X05_Y0E_lo_out[6:5],Tile_X05_Y0E_hi_out[5],Tile_X05_Y0E_lo_out[4],Tile_X05_Y0E_hi_out[4],Tile_X05_Y0E_lo_out[3],Tile_X05_Y0E_lo_out[3:2],Tile_X05_Y0E_lo_out[2],Tile_X05_Y0E_hi_out[2:1],Tile_X05_Y0E_hi_out[1],Tile_X05_Y0E_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X05_Y0E_tile_id (
    .in(Tile_X05_Y0E_tile_id_in),
    .out(Tile_X05_Y0E_tile_id_out)
);
Tile_PE Tile_X05_Y0F (
    .SB_T0_EAST_SB_IN_B1(Tile_X06_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X06_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X05_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X05_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X05_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X05_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X05_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X05_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X05_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X05_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X05_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X05_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X04_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X04_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X05_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X05_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X06_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X06_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X05_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X05_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X05_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X05_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X05_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X05_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X05_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X05_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X05_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X05_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X04_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X04_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X05_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X05_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X06_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X06_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X05_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X05_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X05_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X05_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X05_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X05_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X05_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X05_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X05_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X05_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X04_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X04_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X05_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X05_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X06_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X06_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X05_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X05_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X05_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X05_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X05_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X05_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X05_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X05_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X05_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X05_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X04_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X04_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X05_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X05_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X06_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X06_Y0F_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X05_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X05_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X05_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X05_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X05_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X05_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X05_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X05_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X05_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X05_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X04_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X04_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X05_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X05_Y0F_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X05_Y0E_clk_out),
    .clk_out(Tile_X05_Y0F_clk_out),
    .clk_pass_through(Tile_X05_Y0E_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X05_Y0F_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X05_Y0F_clk_pass_through_out_right),
    .config_config_addr(Tile_X05_Y0E_config_out_config_addr),
    .config_config_data(Tile_X05_Y0E_config_out_config_data),
    .config_out_config_addr(Tile_X05_Y0F_config_out_config_addr),
    .config_out_config_data(Tile_X05_Y0F_config_out_config_data),
    .config_out_read(Tile_X05_Y0F_config_out_read),
    .config_out_write(Tile_X05_Y0F_config_out_write),
    .config_read(Tile_X05_Y0E_config_out_read),
    .config_write(Tile_X05_Y0E_config_out_write),
    .hi(Tile_X05_Y0F_hi_unq1),
    .lo(Tile_X05_Y0F_lo_unq1),
    .read_config_data(Tile_X05_Y0F_read_config_data),
    .read_config_data_in(Tile_X05_Y0E_read_config_data),
    .reset(Tile_X05_Y0E_reset_out),
    .reset_out(Tile_X05_Y0F_reset_out),
    .stall(Tile_X05_Y0E_stall_out),
    .stall_out(Tile_X05_Y0F_stall_out),
    .tile_id(Tile_X05_Y0F_tile_id_in)
);
mantle_wire__typeBit9 Tile_X05_Y0F_hi (
    .in(Tile_X05_Y0F_hi_unq1),
    .out(Tile_X05_Y0F_hi_out)
);
mantle_wire__typeBit8 Tile_X05_Y0F_lo (
    .in(Tile_X05_Y0F_lo_unq1),
    .out(Tile_X05_Y0F_lo_out)
);
wire [15:0] Tile_X05_Y0F_tile_id_out;
assign Tile_X05_Y0F_tile_id_out = {Tile_X05_Y0F_lo_out[7],Tile_X05_Y0F_lo_out[7:6],Tile_X05_Y0F_lo_out[6:5],Tile_X05_Y0F_hi_out[5],Tile_X05_Y0F_lo_out[4],Tile_X05_Y0F_hi_out[4],Tile_X05_Y0F_lo_out[3],Tile_X05_Y0F_lo_out[3:2],Tile_X05_Y0F_lo_out[2],Tile_X05_Y0F_hi_out[2:1],Tile_X05_Y0F_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X05_Y0F_tile_id (
    .in(Tile_X05_Y0F_tile_id_in),
    .out(Tile_X05_Y0F_tile_id_out)
);
Tile_PE Tile_X05_Y10 (
    .SB_T0_EAST_SB_IN_B1(Tile_X06_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X06_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X05_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X05_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X05_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X05_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X05_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X05_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T0_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X05_Y10_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X05_Y10_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X04_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X04_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X05_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X05_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X06_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X06_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X05_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X05_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X05_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X05_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X05_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X05_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T1_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X05_Y10_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X05_Y10_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X04_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X04_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X05_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X05_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X06_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X06_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X05_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X05_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X05_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X05_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X05_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X05_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T2_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X05_Y10_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X05_Y10_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X04_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X04_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X05_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X05_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X06_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X06_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X05_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X05_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X05_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X05_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X05_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X05_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T3_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X05_Y10_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X05_Y10_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X04_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X04_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X05_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X05_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X06_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X06_Y10_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X05_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X05_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X05_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X05_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X05_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X05_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T4_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X05_Y10_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X05_Y10_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X04_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X04_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X05_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X05_Y10_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X05_Y0F_clk_out),
    .clk_out(Tile_X05_Y10_clk_out),
    .clk_pass_through(Tile_X05_Y0F_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X05_Y10_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X05_Y10_clk_pass_through_out_right),
    .config_config_addr(Tile_X05_Y0F_config_out_config_addr),
    .config_config_data(Tile_X05_Y0F_config_out_config_data),
    .config_out_config_addr(Tile_X05_Y10_config_out_config_addr),
    .config_out_config_data(Tile_X05_Y10_config_out_config_data),
    .config_out_read(Tile_X05_Y10_config_out_read),
    .config_out_write(Tile_X05_Y10_config_out_write),
    .config_read(Tile_X05_Y0F_config_out_read),
    .config_write(Tile_X05_Y0F_config_out_write),
    .hi(Tile_X05_Y10_hi),
    .lo(Tile_X05_Y10_lo_unq1),
    .read_config_data(Tile_X05_Y10_read_config_data),
    .read_config_data_in(Tile_X05_Y0F_read_config_data),
    .reset(Tile_X05_Y0F_reset_out),
    .reset_out(Tile_X05_Y10_reset_out),
    .stall(Tile_X05_Y0F_stall_out),
    .stall_out(Tile_X05_Y10_stall_out),
    .tile_id(Tile_X05_Y10_tile_id_in)
);
mantle_wire__typeBit8 Tile_X05_Y10_lo (
    .in(Tile_X05_Y10_lo_unq1),
    .out(Tile_X05_Y10_lo_out)
);
wire [15:0] Tile_X05_Y10_tile_id_out;
assign Tile_X05_Y10_tile_id_out = {Tile_X05_Y10_lo_out[7],Tile_X05_Y10_lo_out[7:6],Tile_X05_Y10_lo_out[6:5],Tile_X05_Y10_hi[5],Tile_X05_Y10_lo_out[4],Tile_X05_Y10_hi[4],Tile_X05_Y10_lo_out[3],Tile_X05_Y10_lo_out[3:2],Tile_X05_Y10_hi[2],Tile_X05_Y10_lo_out[1],Tile_X05_Y10_lo_out[1:0],Tile_X05_Y10_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X05_Y10_tile_id (
    .in(Tile_X05_Y10_tile_id_in),
    .out(Tile_X05_Y10_tile_id_out)
);
wire [15:0] Tile_X06_Y00_tile_id;
assign Tile_X06_Y00_tile_id = {Tile_X06_Y00_lo[7],Tile_X06_Y00_lo[7:6],Tile_X06_Y00_lo[6:5],Tile_X06_Y00_hi[5],Tile_X06_Y00_hi[5],Tile_X06_Y00_lo[4:3],Tile_X06_Y00_lo[3:2],Tile_X06_Y00_lo[2:1],Tile_X06_Y00_lo[1:0],Tile_X06_Y00_lo[0]};
Tile_io_core Tile_X06_Y00 (
    .tile_id(Tile_X06_Y00_tile_id),
    .glb2io_1(glb2io_1_X06_Y00),
    .f2io_1(Tile_X06_Y01_SB_T0_NORTH_SB_OUT_B1),
    .io2glb_1(Tile_X06_Y00_io2glb_1),
    .io2f_1(Tile_X06_Y00_io2f_1),
    .glb2io_16(glb2io_16_X06_Y00),
    .f2io_16(Tile_X06_Y01_SB_T0_NORTH_SB_OUT_B16),
    .io2glb_16(Tile_X06_Y00_io2glb_16),
    .io2f_16(Tile_X06_Y00_io2f_16),
    .hi(Tile_X06_Y00_hi),
    .lo(Tile_X06_Y00_lo)
);
Tile_PE Tile_X06_Y01 (
    .SB_T0_EAST_SB_IN_B1(Tile_X07_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X07_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X06_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X06_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X06_Y00_io2f_1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X06_Y00_io2f_16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X06_Y01_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X06_Y01_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X06_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X06_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X06_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X06_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X05_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X05_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X06_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X06_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X07_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X07_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X06_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X06_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X06_Y00_io2f_1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X06_Y00_io2f_16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X06_Y01_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X06_Y01_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X06_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X06_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X06_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X06_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X05_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X05_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X06_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X06_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X07_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X07_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X06_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X06_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X06_Y00_io2f_1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X06_Y00_io2f_16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X06_Y01_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X06_Y01_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X06_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X06_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X06_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X06_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X05_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X05_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X06_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X06_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X07_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X07_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X06_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X06_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X06_Y00_io2f_1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X06_Y00_io2f_16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X06_Y01_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X06_Y01_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X06_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X06_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X06_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X06_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X05_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X05_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X06_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X06_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X07_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X07_Y01_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X06_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X06_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X06_Y00_io2f_1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X06_Y00_io2f_16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X06_Y01_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X06_Y01_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X06_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X06_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X06_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X06_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X05_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X05_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X06_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X06_Y01_SB_T4_WEST_SB_OUT_B16),
    .clk(clk),
    .clk_out(Tile_X06_Y01_clk_out),
    .clk_pass_through(clk),
    .clk_pass_through_out_bot(Tile_X06_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X06_Y01_clk_pass_through_out_right),
    .config_config_addr(config_6_config_addr),
    .config_config_data(config_6_config_data),
    .config_out_config_addr(Tile_X06_Y01_config_out_config_addr),
    .config_out_config_data(Tile_X06_Y01_config_out_config_data),
    .config_out_read(Tile_X06_Y01_config_out_read),
    .config_out_write(Tile_X06_Y01_config_out_write),
    .config_read(config_6_read),
    .config_write(config_6_write),
    .hi(Tile_X06_Y01_hi),
    .lo(Tile_X06_Y01_lo_unq1),
    .read_config_data(Tile_X06_Y01_read_config_data),
    .read_config_data_in(const_0_32_out),
    .reset(reset),
    .reset_out(Tile_X06_Y01_reset_out),
    .stall(stall[6]),
    .stall_out(Tile_X06_Y01_stall_out),
    .tile_id(Tile_X06_Y01_tile_id_in)
);
mantle_wire__typeBit8 Tile_X06_Y01_lo (
    .in(Tile_X06_Y01_lo_unq1),
    .out(Tile_X06_Y01_lo_out)
);
wire [15:0] Tile_X06_Y01_tile_id_out;
assign Tile_X06_Y01_tile_id_out = {Tile_X06_Y01_lo_out[7],Tile_X06_Y01_lo_out[7:6],Tile_X06_Y01_lo_out[6:5],Tile_X06_Y01_hi[5],Tile_X06_Y01_hi[5],Tile_X06_Y01_lo_out[4:3],Tile_X06_Y01_lo_out[3:2],Tile_X06_Y01_lo_out[2:1],Tile_X06_Y01_lo_out[1:0],Tile_X06_Y01_hi[0]};
mantle_wire__typeBitIn16 Tile_X06_Y01_tile_id (
    .in(Tile_X06_Y01_tile_id_in),
    .out(Tile_X06_Y01_tile_id_out)
);
Tile_PE Tile_X06_Y02 (
    .SB_T0_EAST_SB_IN_B1(Tile_X07_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X07_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X06_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X06_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X06_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X06_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X06_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X06_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X06_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X06_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X06_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X06_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X05_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X05_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X06_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X06_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X07_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X07_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X06_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X06_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X06_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X06_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X06_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X06_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X06_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X06_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X06_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X06_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X05_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X05_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X06_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X06_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X07_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X07_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X06_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X06_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X06_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X06_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X06_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X06_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X06_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X06_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X06_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X06_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X05_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X05_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X06_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X06_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X07_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X07_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X06_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X06_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X06_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X06_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X06_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X06_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X06_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X06_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X06_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X06_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X05_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X05_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X06_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X06_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X07_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X07_Y02_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X06_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X06_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X06_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X06_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X06_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X06_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X06_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X06_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X06_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X06_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X05_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X05_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X06_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X06_Y02_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y01_clk_out),
    .clk_out(Tile_X06_Y02_clk_out),
    .clk_pass_through(Tile_X06_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X06_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X06_Y02_clk_pass_through_out_right),
    .config_config_addr(Tile_X06_Y01_config_out_config_addr),
    .config_config_data(Tile_X06_Y01_config_out_config_data),
    .config_out_config_addr(Tile_X06_Y02_config_out_config_addr),
    .config_out_config_data(Tile_X06_Y02_config_out_config_data),
    .config_out_read(Tile_X06_Y02_config_out_read),
    .config_out_write(Tile_X06_Y02_config_out_write),
    .config_read(Tile_X06_Y01_config_out_read),
    .config_write(Tile_X06_Y01_config_out_write),
    .hi(Tile_X06_Y02_hi),
    .lo(Tile_X06_Y02_lo_unq1),
    .read_config_data(Tile_X06_Y02_read_config_data),
    .read_config_data_in(Tile_X06_Y01_read_config_data),
    .reset(Tile_X06_Y01_reset_out),
    .reset_out(Tile_X06_Y02_reset_out),
    .stall(Tile_X06_Y01_stall_out),
    .stall_out(Tile_X06_Y02_stall_out),
    .tile_id(Tile_X06_Y02_tile_id_in)
);
mantle_wire__typeBit8 Tile_X06_Y02_lo (
    .in(Tile_X06_Y02_lo_unq1),
    .out(Tile_X06_Y02_lo_out)
);
wire [15:0] Tile_X06_Y02_tile_id_out;
assign Tile_X06_Y02_tile_id_out = {Tile_X06_Y02_lo_out[7],Tile_X06_Y02_lo_out[7:6],Tile_X06_Y02_lo_out[6:5],Tile_X06_Y02_hi[5],Tile_X06_Y02_hi[5],Tile_X06_Y02_lo_out[4:3],Tile_X06_Y02_lo_out[3:2],Tile_X06_Y02_lo_out[2:1],Tile_X06_Y02_lo_out[1],Tile_X06_Y02_hi[1],Tile_X06_Y02_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X06_Y02_tile_id (
    .in(Tile_X06_Y02_tile_id_in),
    .out(Tile_X06_Y02_tile_id_out)
);
Tile_PE Tile_X06_Y03 (
    .SB_T0_EAST_SB_IN_B1(Tile_X07_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X07_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X06_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X06_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X06_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X06_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X06_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X06_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X06_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X06_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X06_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X06_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X05_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X05_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X06_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X06_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X07_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X07_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X06_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X06_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X06_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X06_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X06_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X06_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X06_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X06_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X06_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X06_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X05_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X05_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X06_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X06_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X07_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X07_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X06_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X06_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X06_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X06_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X06_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X06_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X06_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X06_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X06_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X06_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X05_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X05_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X06_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X06_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X07_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X07_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X06_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X06_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X06_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X06_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X06_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X06_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X06_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X06_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X06_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X06_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X05_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X05_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X06_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X06_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X07_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X07_Y03_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X06_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X06_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X06_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X06_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X06_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X06_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X06_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X06_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X06_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X06_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X05_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X05_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X06_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X06_Y03_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y02_clk_out),
    .clk_out(Tile_X06_Y03_clk_out),
    .clk_pass_through(Tile_X06_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X06_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X06_Y03_clk_pass_through_out_right),
    .config_config_addr(Tile_X06_Y02_config_out_config_addr),
    .config_config_data(Tile_X06_Y02_config_out_config_data),
    .config_out_config_addr(Tile_X06_Y03_config_out_config_addr),
    .config_out_config_data(Tile_X06_Y03_config_out_config_data),
    .config_out_read(Tile_X06_Y03_config_out_read),
    .config_out_write(Tile_X06_Y03_config_out_write),
    .config_read(Tile_X06_Y02_config_out_read),
    .config_write(Tile_X06_Y02_config_out_write),
    .hi(Tile_X06_Y03_hi_unq1),
    .lo(Tile_X06_Y03_lo_unq1),
    .read_config_data(Tile_X06_Y03_read_config_data),
    .read_config_data_in(Tile_X06_Y02_read_config_data),
    .reset(Tile_X06_Y02_reset_out),
    .reset_out(Tile_X06_Y03_reset_out),
    .stall(Tile_X06_Y02_stall_out),
    .stall_out(Tile_X06_Y03_stall_out),
    .tile_id(Tile_X06_Y03_tile_id_in)
);
mantle_wire__typeBit9 Tile_X06_Y03_hi (
    .in(Tile_X06_Y03_hi_unq1),
    .out(Tile_X06_Y03_hi_out)
);
mantle_wire__typeBit8 Tile_X06_Y03_lo (
    .in(Tile_X06_Y03_lo_unq1),
    .out(Tile_X06_Y03_lo_out)
);
wire [15:0] Tile_X06_Y03_tile_id_out;
assign Tile_X06_Y03_tile_id_out = {Tile_X06_Y03_lo_out[7],Tile_X06_Y03_lo_out[7:6],Tile_X06_Y03_lo_out[6:5],Tile_X06_Y03_hi_out[5],Tile_X06_Y03_hi_out[5],Tile_X06_Y03_lo_out[4:3],Tile_X06_Y03_lo_out[3:2],Tile_X06_Y03_lo_out[2:1],Tile_X06_Y03_lo_out[1],Tile_X06_Y03_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X06_Y03_tile_id (
    .in(Tile_X06_Y03_tile_id_in),
    .out(Tile_X06_Y03_tile_id_out)
);
Tile_PE Tile_X06_Y04 (
    .SB_T0_EAST_SB_IN_B1(Tile_X07_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X07_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X06_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X06_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X06_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X06_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X06_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X06_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X06_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X06_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X06_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X06_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X05_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X05_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X06_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X06_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X07_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X07_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X06_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X06_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X06_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X06_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X06_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X06_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X06_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X06_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X06_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X06_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X05_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X05_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X06_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X06_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X07_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X07_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X06_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X06_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X06_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X06_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X06_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X06_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X06_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X06_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X06_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X06_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X05_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X05_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X06_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X06_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X07_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X07_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X06_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X06_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X06_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X06_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X06_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X06_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X06_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X06_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X06_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X06_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X05_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X05_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X06_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X06_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X07_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X07_Y04_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X06_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X06_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X06_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X06_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X06_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X06_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X06_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X06_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X06_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X06_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X05_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X05_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X06_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X06_Y04_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y03_clk_out),
    .clk_out(Tile_X06_Y04_clk_out),
    .clk_pass_through(Tile_X06_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X06_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X06_Y04_clk_pass_through_out_right),
    .config_config_addr(Tile_X06_Y03_config_out_config_addr),
    .config_config_data(Tile_X06_Y03_config_out_config_data),
    .config_out_config_addr(Tile_X06_Y04_config_out_config_addr),
    .config_out_config_data(Tile_X06_Y04_config_out_config_data),
    .config_out_read(Tile_X06_Y04_config_out_read),
    .config_out_write(Tile_X06_Y04_config_out_write),
    .config_read(Tile_X06_Y03_config_out_read),
    .config_write(Tile_X06_Y03_config_out_write),
    .hi(Tile_X06_Y04_hi),
    .lo(Tile_X06_Y04_lo_unq1),
    .read_config_data(Tile_X06_Y04_read_config_data),
    .read_config_data_in(Tile_X06_Y03_read_config_data),
    .reset(Tile_X06_Y03_reset_out),
    .reset_out(Tile_X06_Y04_reset_out),
    .stall(Tile_X06_Y03_stall_out),
    .stall_out(Tile_X06_Y04_stall_out),
    .tile_id(Tile_X06_Y04_tile_id_in)
);
mantle_wire__typeBit8 Tile_X06_Y04_lo (
    .in(Tile_X06_Y04_lo_unq1),
    .out(Tile_X06_Y04_lo_out)
);
wire [15:0] Tile_X06_Y04_tile_id_out;
assign Tile_X06_Y04_tile_id_out = {Tile_X06_Y04_lo_out[7],Tile_X06_Y04_lo_out[7:6],Tile_X06_Y04_lo_out[6:5],Tile_X06_Y04_hi[5],Tile_X06_Y04_hi[5],Tile_X06_Y04_lo_out[4:3],Tile_X06_Y04_lo_out[3:2],Tile_X06_Y04_lo_out[2:1],Tile_X06_Y04_hi[1],Tile_X06_Y04_lo_out[0],Tile_X06_Y04_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X06_Y04_tile_id (
    .in(Tile_X06_Y04_tile_id_in),
    .out(Tile_X06_Y04_tile_id_out)
);
Tile_PE Tile_X06_Y05 (
    .SB_T0_EAST_SB_IN_B1(Tile_X07_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X07_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X06_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X06_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X06_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X06_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X06_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X06_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X06_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X06_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X06_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X06_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X05_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X05_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X06_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X06_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X07_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X07_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X06_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X06_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X06_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X06_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X06_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X06_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X06_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X06_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X06_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X06_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X05_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X05_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X06_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X06_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X07_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X07_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X06_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X06_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X06_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X06_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X06_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X06_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X06_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X06_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X06_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X06_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X05_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X05_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X06_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X06_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X07_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X07_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X06_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X06_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X06_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X06_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X06_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X06_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X06_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X06_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X06_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X06_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X05_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X05_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X06_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X06_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X07_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X07_Y05_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X06_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X06_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X06_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X06_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X06_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X06_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X06_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X06_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X06_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X06_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X05_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X05_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X06_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X06_Y05_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y04_clk_out),
    .clk_out(Tile_X06_Y05_clk_out),
    .clk_pass_through(Tile_X06_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X06_Y05_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X06_Y05_clk_pass_through_out_right),
    .config_config_addr(Tile_X06_Y04_config_out_config_addr),
    .config_config_data(Tile_X06_Y04_config_out_config_data),
    .config_out_config_addr(Tile_X06_Y05_config_out_config_addr),
    .config_out_config_data(Tile_X06_Y05_config_out_config_data),
    .config_out_read(Tile_X06_Y05_config_out_read),
    .config_out_write(Tile_X06_Y05_config_out_write),
    .config_read(Tile_X06_Y04_config_out_read),
    .config_write(Tile_X06_Y04_config_out_write),
    .hi(Tile_X06_Y05_hi),
    .lo(Tile_X06_Y05_lo_unq1),
    .read_config_data(Tile_X06_Y05_read_config_data),
    .read_config_data_in(Tile_X06_Y04_read_config_data),
    .reset(Tile_X06_Y04_reset_out),
    .reset_out(Tile_X06_Y05_reset_out),
    .stall(Tile_X06_Y04_stall_out),
    .stall_out(Tile_X06_Y05_stall_out),
    .tile_id(Tile_X06_Y05_tile_id_in)
);
mantle_wire__typeBit8 Tile_X06_Y05_lo (
    .in(Tile_X06_Y05_lo_unq1),
    .out(Tile_X06_Y05_lo_out)
);
wire [15:0] Tile_X06_Y05_tile_id_out;
assign Tile_X06_Y05_tile_id_out = {Tile_X06_Y05_lo_out[7],Tile_X06_Y05_lo_out[7:6],Tile_X06_Y05_lo_out[6:5],Tile_X06_Y05_hi[5],Tile_X06_Y05_hi[5],Tile_X06_Y05_lo_out[4:3],Tile_X06_Y05_lo_out[3:2],Tile_X06_Y05_lo_out[2:1],Tile_X06_Y05_hi[1],Tile_X06_Y05_lo_out[0],Tile_X06_Y05_hi[0]};
mantle_wire__typeBitIn16 Tile_X06_Y05_tile_id (
    .in(Tile_X06_Y05_tile_id_in),
    .out(Tile_X06_Y05_tile_id_out)
);
Tile_PE Tile_X06_Y06 (
    .SB_T0_EAST_SB_IN_B1(Tile_X07_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X07_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X06_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X06_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X06_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X06_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X06_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X06_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X06_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X06_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X06_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X06_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X05_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X05_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X06_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X06_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X07_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X07_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X06_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X06_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X06_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X06_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X06_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X06_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X06_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X06_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X06_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X06_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X05_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X05_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X06_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X06_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X07_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X07_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X06_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X06_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X06_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X06_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X06_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X06_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X06_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X06_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X06_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X06_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X05_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X05_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X06_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X06_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X07_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X07_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X06_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X06_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X06_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X06_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X06_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X06_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X06_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X06_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X06_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X06_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X05_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X05_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X06_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X06_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X07_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X07_Y06_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X06_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X06_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X06_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X06_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X06_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X06_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X06_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X06_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X06_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X06_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X05_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X05_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X06_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X06_Y06_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y05_clk_out),
    .clk_out(Tile_X06_Y06_clk_out),
    .clk_pass_through(Tile_X06_Y05_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X06_Y06_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X06_Y06_clk_pass_through_out_right),
    .config_config_addr(Tile_X06_Y05_config_out_config_addr),
    .config_config_data(Tile_X06_Y05_config_out_config_data),
    .config_out_config_addr(Tile_X06_Y06_config_out_config_addr),
    .config_out_config_data(Tile_X06_Y06_config_out_config_data),
    .config_out_read(Tile_X06_Y06_config_out_read),
    .config_out_write(Tile_X06_Y06_config_out_write),
    .config_read(Tile_X06_Y05_config_out_read),
    .config_write(Tile_X06_Y05_config_out_write),
    .hi(Tile_X06_Y06_hi),
    .lo(Tile_X06_Y06_lo_unq1),
    .read_config_data(Tile_X06_Y06_read_config_data),
    .read_config_data_in(Tile_X06_Y05_read_config_data),
    .reset(Tile_X06_Y05_reset_out),
    .reset_out(Tile_X06_Y06_reset_out),
    .stall(Tile_X06_Y05_stall_out),
    .stall_out(Tile_X06_Y06_stall_out),
    .tile_id(Tile_X06_Y06_tile_id_in)
);
mantle_wire__typeBit8 Tile_X06_Y06_lo (
    .in(Tile_X06_Y06_lo_unq1),
    .out(Tile_X06_Y06_lo_out)
);
wire [15:0] Tile_X06_Y06_tile_id_out;
assign Tile_X06_Y06_tile_id_out = {Tile_X06_Y06_lo_out[7],Tile_X06_Y06_lo_out[7:6],Tile_X06_Y06_lo_out[6:5],Tile_X06_Y06_hi[5],Tile_X06_Y06_hi[5],Tile_X06_Y06_lo_out[4:3],Tile_X06_Y06_lo_out[3:2],Tile_X06_Y06_lo_out[2:1],Tile_X06_Y06_hi[1],Tile_X06_Y06_hi[1],Tile_X06_Y06_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X06_Y06_tile_id (
    .in(Tile_X06_Y06_tile_id_in),
    .out(Tile_X06_Y06_tile_id_out)
);
Tile_PE Tile_X06_Y07 (
    .SB_T0_EAST_SB_IN_B1(Tile_X07_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X07_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X06_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X06_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X06_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X06_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X06_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X06_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X06_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X06_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X06_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X06_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X05_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X05_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X06_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X06_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X07_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X07_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X06_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X06_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X06_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X06_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X06_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X06_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X06_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X06_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X06_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X06_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X05_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X05_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X06_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X06_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X07_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X07_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X06_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X06_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X06_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X06_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X06_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X06_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X06_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X06_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X06_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X06_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X05_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X05_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X06_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X06_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X07_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X07_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X06_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X06_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X06_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X06_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X06_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X06_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X06_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X06_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X06_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X06_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X05_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X05_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X06_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X06_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X07_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X07_Y07_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X06_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X06_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X06_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X06_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X06_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X06_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X06_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X06_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X06_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X06_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X05_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X05_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X06_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X06_Y07_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y06_clk_out),
    .clk_out(Tile_X06_Y07_clk_out),
    .clk_pass_through(Tile_X06_Y06_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X06_Y07_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X06_Y07_clk_pass_through_out_right),
    .config_config_addr(Tile_X06_Y06_config_out_config_addr),
    .config_config_data(Tile_X06_Y06_config_out_config_data),
    .config_out_config_addr(Tile_X06_Y07_config_out_config_addr),
    .config_out_config_data(Tile_X06_Y07_config_out_config_data),
    .config_out_read(Tile_X06_Y07_config_out_read),
    .config_out_write(Tile_X06_Y07_config_out_write),
    .config_read(Tile_X06_Y06_config_out_read),
    .config_write(Tile_X06_Y06_config_out_write),
    .hi(Tile_X06_Y07_hi_unq1),
    .lo(Tile_X06_Y07_lo_unq1),
    .read_config_data(Tile_X06_Y07_read_config_data),
    .read_config_data_in(Tile_X06_Y06_read_config_data),
    .reset(Tile_X06_Y06_reset_out),
    .reset_out(Tile_X06_Y07_reset_out),
    .stall(Tile_X06_Y06_stall_out),
    .stall_out(Tile_X06_Y07_stall_out),
    .tile_id(Tile_X06_Y07_tile_id_in)
);
mantle_wire__typeBit9 Tile_X06_Y07_hi (
    .in(Tile_X06_Y07_hi_unq1),
    .out(Tile_X06_Y07_hi_out)
);
mantle_wire__typeBit8 Tile_X06_Y07_lo (
    .in(Tile_X06_Y07_lo_unq1),
    .out(Tile_X06_Y07_lo_out)
);
wire [15:0] Tile_X06_Y07_tile_id_out;
assign Tile_X06_Y07_tile_id_out = {Tile_X06_Y07_lo_out[7],Tile_X06_Y07_lo_out[7:6],Tile_X06_Y07_lo_out[6:5],Tile_X06_Y07_hi_out[5],Tile_X06_Y07_hi_out[5],Tile_X06_Y07_lo_out[4:3],Tile_X06_Y07_lo_out[3:2],Tile_X06_Y07_lo_out[2:1],Tile_X06_Y07_hi_out[1],Tile_X06_Y07_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X06_Y07_tile_id (
    .in(Tile_X06_Y07_tile_id_in),
    .out(Tile_X06_Y07_tile_id_out)
);
Tile_PE Tile_X06_Y08 (
    .SB_T0_EAST_SB_IN_B1(Tile_X07_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X07_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X06_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X06_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X06_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X06_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X06_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X06_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X06_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X06_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X06_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X06_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X05_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X05_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X06_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X06_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X07_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X07_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X06_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X06_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X06_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X06_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X06_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X06_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X06_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X06_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X06_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X06_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X05_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X05_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X06_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X06_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X07_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X07_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X06_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X06_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X06_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X06_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X06_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X06_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X06_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X06_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X06_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X06_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X05_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X05_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X06_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X06_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X07_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X07_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X06_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X06_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X06_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X06_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X06_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X06_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X06_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X06_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X06_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X06_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X05_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X05_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X06_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X06_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X07_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X07_Y08_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X06_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X06_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X06_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X06_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X06_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X06_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X06_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X06_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X06_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X06_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X05_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X05_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X06_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X06_Y08_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y07_clk_out),
    .clk_out(Tile_X06_Y08_clk_out),
    .clk_pass_through(Tile_X06_Y07_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X06_Y08_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X06_Y08_clk_pass_through_out_right),
    .config_config_addr(Tile_X06_Y07_config_out_config_addr),
    .config_config_data(Tile_X06_Y07_config_out_config_data),
    .config_out_config_addr(Tile_X06_Y08_config_out_config_addr),
    .config_out_config_data(Tile_X06_Y08_config_out_config_data),
    .config_out_read(Tile_X06_Y08_config_out_read),
    .config_out_write(Tile_X06_Y08_config_out_write),
    .config_read(Tile_X06_Y07_config_out_read),
    .config_write(Tile_X06_Y07_config_out_write),
    .hi(Tile_X06_Y08_hi),
    .lo(Tile_X06_Y08_lo_unq1),
    .read_config_data(Tile_X06_Y08_read_config_data),
    .read_config_data_in(Tile_X06_Y07_read_config_data),
    .reset(Tile_X06_Y07_reset_out),
    .reset_out(Tile_X06_Y08_reset_out),
    .stall(Tile_X06_Y07_stall_out),
    .stall_out(Tile_X06_Y08_stall_out),
    .tile_id(Tile_X06_Y08_tile_id_in)
);
mantle_wire__typeBit8 Tile_X06_Y08_lo (
    .in(Tile_X06_Y08_lo_unq1),
    .out(Tile_X06_Y08_lo_out)
);
wire [15:0] Tile_X06_Y08_tile_id_out;
assign Tile_X06_Y08_tile_id_out = {Tile_X06_Y08_lo_out[7],Tile_X06_Y08_lo_out[7:6],Tile_X06_Y08_lo_out[6:5],Tile_X06_Y08_hi[5],Tile_X06_Y08_hi[5],Tile_X06_Y08_lo_out[4:3],Tile_X06_Y08_lo_out[3:2],Tile_X06_Y08_lo_out[2],Tile_X06_Y08_hi[2],Tile_X06_Y08_lo_out[1:0],Tile_X06_Y08_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X06_Y08_tile_id (
    .in(Tile_X06_Y08_tile_id_in),
    .out(Tile_X06_Y08_tile_id_out)
);
Tile_PE Tile_X06_Y09 (
    .SB_T0_EAST_SB_IN_B1(Tile_X07_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X07_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X06_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X06_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X06_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X06_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X06_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X06_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X06_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X06_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X06_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X06_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X05_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X05_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X06_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X06_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X07_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X07_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X06_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X06_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X06_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X06_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X06_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X06_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X06_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X06_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X06_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X06_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X05_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X05_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X06_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X06_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X07_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X07_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X06_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X06_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X06_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X06_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X06_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X06_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X06_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X06_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X06_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X06_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X05_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X05_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X06_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X06_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X07_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X07_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X06_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X06_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X06_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X06_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X06_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X06_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X06_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X06_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X06_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X06_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X05_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X05_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X06_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X06_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X07_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X07_Y09_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X06_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X06_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X06_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X06_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X06_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X06_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X06_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X06_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X06_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X06_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X05_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X05_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X06_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X06_Y09_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y08_clk_out),
    .clk_out(Tile_X06_Y09_clk_out),
    .clk_pass_through(Tile_X06_Y08_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X06_Y09_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X06_Y09_clk_pass_through_out_right),
    .config_config_addr(ConfigPipeStage_inst6_config_out_config_addr),
    .config_config_data(ConfigPipeStage_inst6_config_out_config_data),
    .config_out_config_addr(Tile_X06_Y09_config_out_config_addr),
    .config_out_config_data(Tile_X06_Y09_config_out_config_data),
    .config_out_read(Tile_X06_Y09_config_out_read),
    .config_out_write(Tile_X06_Y09_config_out_write),
    .config_read(ConfigPipeStage_inst6_config_out_read),
    .config_write(ConfigPipeStage_inst6_config_out_write),
    .hi(Tile_X06_Y09_hi),
    .lo(Tile_X06_Y09_lo_unq1),
    .read_config_data(Tile_X06_Y09_read_config_data),
    .read_config_data_in(Tile_X06_Y08_read_config_data),
    .reset(Tile_X06_Y08_reset_out),
    .reset_out(Tile_X06_Y09_reset_out),
    .stall(Tile_X06_Y08_stall_out),
    .stall_out(Tile_X06_Y09_stall_out),
    .tile_id(Tile_X06_Y09_tile_id_in)
);
mantle_wire__typeBit8 Tile_X06_Y09_lo (
    .in(Tile_X06_Y09_lo_unq1),
    .out(Tile_X06_Y09_lo_out)
);
wire [15:0] Tile_X06_Y09_tile_id_out;
assign Tile_X06_Y09_tile_id_out = {Tile_X06_Y09_lo_out[7],Tile_X06_Y09_lo_out[7:6],Tile_X06_Y09_lo_out[6:5],Tile_X06_Y09_hi[5],Tile_X06_Y09_hi[5],Tile_X06_Y09_lo_out[4:3],Tile_X06_Y09_lo_out[3:2],Tile_X06_Y09_lo_out[2],Tile_X06_Y09_hi[2],Tile_X06_Y09_lo_out[1:0],Tile_X06_Y09_hi[0]};
mantle_wire__typeBitIn16 Tile_X06_Y09_tile_id (
    .in(Tile_X06_Y09_tile_id_in),
    .out(Tile_X06_Y09_tile_id_out)
);
Tile_PE Tile_X06_Y0A (
    .SB_T0_EAST_SB_IN_B1(Tile_X07_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X07_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X06_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X06_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X06_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X06_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X06_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X06_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X06_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X06_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X06_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X06_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X05_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X05_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X06_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X06_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X07_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X07_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X06_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X06_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X06_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X06_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X06_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X06_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X06_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X06_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X06_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X06_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X05_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X05_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X06_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X06_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X07_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X07_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X06_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X06_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X06_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X06_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X06_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X06_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X06_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X06_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X06_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X06_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X05_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X05_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X06_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X06_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X07_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X07_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X06_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X06_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X06_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X06_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X06_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X06_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X06_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X06_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X06_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X06_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X05_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X05_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X06_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X06_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X07_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X07_Y0A_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X06_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X06_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X06_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X06_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X06_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X06_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X06_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X06_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X06_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X06_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X05_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X05_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X06_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X06_Y0A_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y09_clk_out),
    .clk_out(Tile_X06_Y0A_clk_out),
    .clk_pass_through(Tile_X06_Y09_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X06_Y0A_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X06_Y0A_clk_pass_through_out_right),
    .config_config_addr(Tile_X06_Y09_config_out_config_addr),
    .config_config_data(Tile_X06_Y09_config_out_config_data),
    .config_out_config_addr(Tile_X06_Y0A_config_out_config_addr),
    .config_out_config_data(Tile_X06_Y0A_config_out_config_data),
    .config_out_read(Tile_X06_Y0A_config_out_read),
    .config_out_write(Tile_X06_Y0A_config_out_write),
    .config_read(Tile_X06_Y09_config_out_read),
    .config_write(Tile_X06_Y09_config_out_write),
    .hi(Tile_X06_Y0A_hi),
    .lo(Tile_X06_Y0A_lo_unq1),
    .read_config_data(Tile_X06_Y0A_read_config_data),
    .read_config_data_in(Tile_X06_Y09_read_config_data),
    .reset(Tile_X06_Y09_reset_out),
    .reset_out(Tile_X06_Y0A_reset_out),
    .stall(Tile_X06_Y09_stall_out),
    .stall_out(Tile_X06_Y0A_stall_out),
    .tile_id(Tile_X06_Y0A_tile_id_in)
);
mantle_wire__typeBit8 Tile_X06_Y0A_lo (
    .in(Tile_X06_Y0A_lo_unq1),
    .out(Tile_X06_Y0A_lo_out)
);
wire [15:0] Tile_X06_Y0A_tile_id_out;
assign Tile_X06_Y0A_tile_id_out = {Tile_X06_Y0A_lo_out[7],Tile_X06_Y0A_lo_out[7:6],Tile_X06_Y0A_lo_out[6:5],Tile_X06_Y0A_hi[5],Tile_X06_Y0A_hi[5],Tile_X06_Y0A_lo_out[4:3],Tile_X06_Y0A_lo_out[3:2],Tile_X06_Y0A_lo_out[2],Tile_X06_Y0A_hi[2],Tile_X06_Y0A_lo_out[1],Tile_X06_Y0A_hi[1],Tile_X06_Y0A_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X06_Y0A_tile_id (
    .in(Tile_X06_Y0A_tile_id_in),
    .out(Tile_X06_Y0A_tile_id_out)
);
Tile_PE Tile_X06_Y0B (
    .SB_T0_EAST_SB_IN_B1(Tile_X07_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X07_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X06_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X06_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X06_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X06_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X06_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X06_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X06_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X06_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X06_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X06_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X05_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X05_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X06_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X06_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X07_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X07_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X06_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X06_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X06_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X06_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X06_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X06_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X06_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X06_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X06_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X06_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X05_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X05_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X06_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X06_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X07_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X07_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X06_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X06_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X06_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X06_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X06_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X06_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X06_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X06_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X06_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X06_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X05_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X05_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X06_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X06_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X07_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X07_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X06_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X06_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X06_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X06_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X06_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X06_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X06_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X06_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X06_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X06_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X05_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X05_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X06_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X06_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X07_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X07_Y0B_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X06_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X06_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X06_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X06_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X06_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X06_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X06_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X06_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X06_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X06_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X05_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X05_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X06_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X06_Y0B_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y0A_clk_out),
    .clk_out(Tile_X06_Y0B_clk_out),
    .clk_pass_through(Tile_X06_Y0A_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X06_Y0B_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X06_Y0B_clk_pass_through_out_right),
    .config_config_addr(Tile_X06_Y0A_config_out_config_addr),
    .config_config_data(Tile_X06_Y0A_config_out_config_data),
    .config_out_config_addr(Tile_X06_Y0B_config_out_config_addr),
    .config_out_config_data(Tile_X06_Y0B_config_out_config_data),
    .config_out_read(Tile_X06_Y0B_config_out_read),
    .config_out_write(Tile_X06_Y0B_config_out_write),
    .config_read(Tile_X06_Y0A_config_out_read),
    .config_write(Tile_X06_Y0A_config_out_write),
    .hi(Tile_X06_Y0B_hi_unq1),
    .lo(Tile_X06_Y0B_lo_unq1),
    .read_config_data(Tile_X06_Y0B_read_config_data),
    .read_config_data_in(Tile_X06_Y0A_read_config_data),
    .reset(Tile_X06_Y0A_reset_out),
    .reset_out(Tile_X06_Y0B_reset_out),
    .stall(Tile_X06_Y0A_stall_out),
    .stall_out(Tile_X06_Y0B_stall_out),
    .tile_id(Tile_X06_Y0B_tile_id_in)
);
mantle_wire__typeBit9 Tile_X06_Y0B_hi (
    .in(Tile_X06_Y0B_hi_unq1),
    .out(Tile_X06_Y0B_hi_out)
);
mantle_wire__typeBit8 Tile_X06_Y0B_lo (
    .in(Tile_X06_Y0B_lo_unq1),
    .out(Tile_X06_Y0B_lo_out)
);
wire [15:0] Tile_X06_Y0B_tile_id_out;
assign Tile_X06_Y0B_tile_id_out = {Tile_X06_Y0B_lo_out[7],Tile_X06_Y0B_lo_out[7:6],Tile_X06_Y0B_lo_out[6:5],Tile_X06_Y0B_hi_out[5],Tile_X06_Y0B_hi_out[5],Tile_X06_Y0B_lo_out[4:3],Tile_X06_Y0B_lo_out[3:2],Tile_X06_Y0B_lo_out[2],Tile_X06_Y0B_hi_out[2],Tile_X06_Y0B_lo_out[1],Tile_X06_Y0B_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X06_Y0B_tile_id (
    .in(Tile_X06_Y0B_tile_id_in),
    .out(Tile_X06_Y0B_tile_id_out)
);
Tile_PE Tile_X06_Y0C (
    .SB_T0_EAST_SB_IN_B1(Tile_X07_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X07_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X06_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X06_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X06_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X06_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X06_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X06_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X06_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X06_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X06_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X06_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X05_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X05_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X06_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X06_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X07_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X07_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X06_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X06_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X06_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X06_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X06_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X06_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X06_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X06_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X06_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X06_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X05_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X05_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X06_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X06_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X07_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X07_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X06_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X06_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X06_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X06_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X06_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X06_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X06_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X06_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X06_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X06_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X05_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X05_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X06_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X06_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X07_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X07_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X06_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X06_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X06_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X06_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X06_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X06_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X06_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X06_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X06_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X06_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X05_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X05_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X06_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X06_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X07_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X07_Y0C_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X06_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X06_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X06_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X06_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X06_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X06_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X06_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X06_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X06_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X06_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X05_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X05_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X06_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X06_Y0C_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y0B_clk_out),
    .clk_out(Tile_X06_Y0C_clk_out),
    .clk_pass_through(Tile_X06_Y0B_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X06_Y0C_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X06_Y0C_clk_pass_through_out_right),
    .config_config_addr(Tile_X06_Y0B_config_out_config_addr),
    .config_config_data(Tile_X06_Y0B_config_out_config_data),
    .config_out_config_addr(Tile_X06_Y0C_config_out_config_addr),
    .config_out_config_data(Tile_X06_Y0C_config_out_config_data),
    .config_out_read(Tile_X06_Y0C_config_out_read),
    .config_out_write(Tile_X06_Y0C_config_out_write),
    .config_read(Tile_X06_Y0B_config_out_read),
    .config_write(Tile_X06_Y0B_config_out_write),
    .hi(Tile_X06_Y0C_hi_unq1),
    .lo(Tile_X06_Y0C_lo_unq1),
    .read_config_data(Tile_X06_Y0C_read_config_data),
    .read_config_data_in(Tile_X06_Y0B_read_config_data),
    .reset(Tile_X06_Y0B_reset_out),
    .reset_out(Tile_X06_Y0C_reset_out),
    .stall(Tile_X06_Y0B_stall_out),
    .stall_out(Tile_X06_Y0C_stall_out),
    .tile_id(Tile_X06_Y0C_tile_id_in)
);
mantle_wire__typeBit9 Tile_X06_Y0C_hi (
    .in(Tile_X06_Y0C_hi_unq1),
    .out(Tile_X06_Y0C_hi_out)
);
mantle_wire__typeBit8 Tile_X06_Y0C_lo (
    .in(Tile_X06_Y0C_lo_unq1),
    .out(Tile_X06_Y0C_lo_out)
);
wire [15:0] Tile_X06_Y0C_tile_id_out;
assign Tile_X06_Y0C_tile_id_out = {Tile_X06_Y0C_lo_out[7],Tile_X06_Y0C_lo_out[7:6],Tile_X06_Y0C_lo_out[6:5],Tile_X06_Y0C_hi_out[5],Tile_X06_Y0C_hi_out[5],Tile_X06_Y0C_lo_out[4:3],Tile_X06_Y0C_lo_out[3:2],Tile_X06_Y0C_lo_out[2],Tile_X06_Y0C_hi_out[2:1],Tile_X06_Y0C_lo_out[0],Tile_X06_Y0C_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X06_Y0C_tile_id (
    .in(Tile_X06_Y0C_tile_id_in),
    .out(Tile_X06_Y0C_tile_id_out)
);
Tile_PE Tile_X06_Y0D (
    .SB_T0_EAST_SB_IN_B1(Tile_X07_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X07_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X06_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X06_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X06_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X06_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X06_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X06_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X06_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X06_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X06_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X06_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X05_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X05_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X06_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X06_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X07_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X07_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X06_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X06_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X06_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X06_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X06_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X06_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X06_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X06_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X06_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X06_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X05_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X05_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X06_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X06_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X07_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X07_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X06_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X06_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X06_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X06_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X06_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X06_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X06_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X06_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X06_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X06_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X05_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X05_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X06_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X06_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X07_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X07_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X06_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X06_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X06_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X06_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X06_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X06_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X06_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X06_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X06_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X06_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X05_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X05_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X06_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X06_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X07_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X07_Y0D_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X06_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X06_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X06_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X06_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X06_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X06_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X06_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X06_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X06_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X06_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X05_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X05_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X06_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X06_Y0D_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y0C_clk_out),
    .clk_out(Tile_X06_Y0D_clk_out),
    .clk_pass_through(Tile_X06_Y0C_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X06_Y0D_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X06_Y0D_clk_pass_through_out_right),
    .config_config_addr(Tile_X06_Y0C_config_out_config_addr),
    .config_config_data(Tile_X06_Y0C_config_out_config_data),
    .config_out_config_addr(Tile_X06_Y0D_config_out_config_addr),
    .config_out_config_data(Tile_X06_Y0D_config_out_config_data),
    .config_out_read(Tile_X06_Y0D_config_out_read),
    .config_out_write(Tile_X06_Y0D_config_out_write),
    .config_read(Tile_X06_Y0C_config_out_read),
    .config_write(Tile_X06_Y0C_config_out_write),
    .hi(Tile_X06_Y0D_hi_unq1),
    .lo(Tile_X06_Y0D_lo_unq1),
    .read_config_data(Tile_X06_Y0D_read_config_data),
    .read_config_data_in(Tile_X06_Y0C_read_config_data),
    .reset(Tile_X06_Y0C_reset_out),
    .reset_out(Tile_X06_Y0D_reset_out),
    .stall(Tile_X06_Y0C_stall_out),
    .stall_out(Tile_X06_Y0D_stall_out),
    .tile_id(Tile_X06_Y0D_tile_id_in)
);
mantle_wire__typeBit9 Tile_X06_Y0D_hi (
    .in(Tile_X06_Y0D_hi_unq1),
    .out(Tile_X06_Y0D_hi_out)
);
mantle_wire__typeBit8 Tile_X06_Y0D_lo (
    .in(Tile_X06_Y0D_lo_unq1),
    .out(Tile_X06_Y0D_lo_out)
);
wire [15:0] Tile_X06_Y0D_tile_id_out;
assign Tile_X06_Y0D_tile_id_out = {Tile_X06_Y0D_lo_out[7],Tile_X06_Y0D_lo_out[7:6],Tile_X06_Y0D_lo_out[6:5],Tile_X06_Y0D_hi_out[5],Tile_X06_Y0D_hi_out[5],Tile_X06_Y0D_lo_out[4:3],Tile_X06_Y0D_lo_out[3:2],Tile_X06_Y0D_lo_out[2],Tile_X06_Y0D_hi_out[2:1],Tile_X06_Y0D_lo_out[0],Tile_X06_Y0D_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X06_Y0D_tile_id (
    .in(Tile_X06_Y0D_tile_id_in),
    .out(Tile_X06_Y0D_tile_id_out)
);
Tile_PE Tile_X06_Y0E (
    .SB_T0_EAST_SB_IN_B1(Tile_X07_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X07_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X06_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X06_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X06_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X06_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X06_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X06_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X06_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X06_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X06_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X06_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X05_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X05_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X06_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X06_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X07_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X07_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X06_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X06_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X06_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X06_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X06_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X06_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X06_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X06_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X06_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X06_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X05_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X05_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X06_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X06_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X07_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X07_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X06_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X06_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X06_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X06_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X06_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X06_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X06_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X06_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X06_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X06_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X05_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X05_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X06_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X06_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X07_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X07_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X06_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X06_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X06_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X06_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X06_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X06_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X06_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X06_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X06_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X06_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X05_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X05_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X06_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X06_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X07_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X07_Y0E_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X06_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X06_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X06_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X06_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X06_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X06_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X06_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X06_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X06_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X06_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X05_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X05_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X06_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X06_Y0E_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y0D_clk_out),
    .clk_out(Tile_X06_Y0E_clk_out),
    .clk_pass_through(Tile_X06_Y0D_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X06_Y0E_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X06_Y0E_clk_pass_through_out_right),
    .config_config_addr(Tile_X06_Y0D_config_out_config_addr),
    .config_config_data(Tile_X06_Y0D_config_out_config_data),
    .config_out_config_addr(Tile_X06_Y0E_config_out_config_addr),
    .config_out_config_data(Tile_X06_Y0E_config_out_config_data),
    .config_out_read(Tile_X06_Y0E_config_out_read),
    .config_out_write(Tile_X06_Y0E_config_out_write),
    .config_read(Tile_X06_Y0D_config_out_read),
    .config_write(Tile_X06_Y0D_config_out_write),
    .hi(Tile_X06_Y0E_hi_unq1),
    .lo(Tile_X06_Y0E_lo_unq1),
    .read_config_data(Tile_X06_Y0E_read_config_data),
    .read_config_data_in(Tile_X06_Y0D_read_config_data),
    .reset(Tile_X06_Y0D_reset_out),
    .reset_out(Tile_X06_Y0E_reset_out),
    .stall(Tile_X06_Y0D_stall_out),
    .stall_out(Tile_X06_Y0E_stall_out),
    .tile_id(Tile_X06_Y0E_tile_id_in)
);
mantle_wire__typeBit9 Tile_X06_Y0E_hi (
    .in(Tile_X06_Y0E_hi_unq1),
    .out(Tile_X06_Y0E_hi_out)
);
mantle_wire__typeBit8 Tile_X06_Y0E_lo (
    .in(Tile_X06_Y0E_lo_unq1),
    .out(Tile_X06_Y0E_lo_out)
);
wire [15:0] Tile_X06_Y0E_tile_id_out;
assign Tile_X06_Y0E_tile_id_out = {Tile_X06_Y0E_lo_out[7],Tile_X06_Y0E_lo_out[7:6],Tile_X06_Y0E_lo_out[6:5],Tile_X06_Y0E_hi_out[5],Tile_X06_Y0E_hi_out[5],Tile_X06_Y0E_lo_out[4:3],Tile_X06_Y0E_lo_out[3:2],Tile_X06_Y0E_lo_out[2],Tile_X06_Y0E_hi_out[2:1],Tile_X06_Y0E_hi_out[1],Tile_X06_Y0E_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X06_Y0E_tile_id (
    .in(Tile_X06_Y0E_tile_id_in),
    .out(Tile_X06_Y0E_tile_id_out)
);
Tile_PE Tile_X06_Y0F (
    .SB_T0_EAST_SB_IN_B1(Tile_X07_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X07_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X06_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X06_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X06_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X06_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X06_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X06_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X06_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X06_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X06_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X06_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X05_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X05_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X06_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X06_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X07_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X07_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X06_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X06_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X06_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X06_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X06_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X06_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X06_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X06_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X06_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X06_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X05_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X05_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X06_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X06_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X07_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X07_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X06_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X06_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X06_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X06_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X06_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X06_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X06_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X06_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X06_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X06_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X05_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X05_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X06_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X06_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X07_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X07_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X06_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X06_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X06_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X06_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X06_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X06_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X06_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X06_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X06_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X06_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X05_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X05_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X06_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X06_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X07_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X07_Y0F_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X06_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X06_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X06_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X06_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X06_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X06_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X06_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X06_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X06_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X06_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X05_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X05_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X06_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X06_Y0F_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y0E_clk_out),
    .clk_out(Tile_X06_Y0F_clk_out),
    .clk_pass_through(Tile_X06_Y0E_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X06_Y0F_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X06_Y0F_clk_pass_through_out_right),
    .config_config_addr(Tile_X06_Y0E_config_out_config_addr),
    .config_config_data(Tile_X06_Y0E_config_out_config_data),
    .config_out_config_addr(Tile_X06_Y0F_config_out_config_addr),
    .config_out_config_data(Tile_X06_Y0F_config_out_config_data),
    .config_out_read(Tile_X06_Y0F_config_out_read),
    .config_out_write(Tile_X06_Y0F_config_out_write),
    .config_read(Tile_X06_Y0E_config_out_read),
    .config_write(Tile_X06_Y0E_config_out_write),
    .hi(Tile_X06_Y0F_hi_unq1),
    .lo(Tile_X06_Y0F_lo_unq1),
    .read_config_data(Tile_X06_Y0F_read_config_data),
    .read_config_data_in(Tile_X06_Y0E_read_config_data),
    .reset(Tile_X06_Y0E_reset_out),
    .reset_out(Tile_X06_Y0F_reset_out),
    .stall(Tile_X06_Y0E_stall_out),
    .stall_out(Tile_X06_Y0F_stall_out),
    .tile_id(Tile_X06_Y0F_tile_id_in)
);
mantle_wire__typeBit9 Tile_X06_Y0F_hi (
    .in(Tile_X06_Y0F_hi_unq1),
    .out(Tile_X06_Y0F_hi_out)
);
mantle_wire__typeBit8 Tile_X06_Y0F_lo (
    .in(Tile_X06_Y0F_lo_unq1),
    .out(Tile_X06_Y0F_lo_out)
);
wire [15:0] Tile_X06_Y0F_tile_id_out;
assign Tile_X06_Y0F_tile_id_out = {Tile_X06_Y0F_lo_out[7],Tile_X06_Y0F_lo_out[7:6],Tile_X06_Y0F_lo_out[6:5],Tile_X06_Y0F_hi_out[5],Tile_X06_Y0F_hi_out[5],Tile_X06_Y0F_lo_out[4:3],Tile_X06_Y0F_lo_out[3:2],Tile_X06_Y0F_lo_out[2],Tile_X06_Y0F_hi_out[2:1],Tile_X06_Y0F_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X06_Y0F_tile_id (
    .in(Tile_X06_Y0F_tile_id_in),
    .out(Tile_X06_Y0F_tile_id_out)
);
Tile_PE Tile_X06_Y10 (
    .SB_T0_EAST_SB_IN_B1(Tile_X07_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X07_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X06_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X06_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X06_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X06_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X06_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X06_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T0_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X06_Y10_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X06_Y10_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X05_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X05_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X06_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X06_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X07_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X07_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X06_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X06_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X06_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X06_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X06_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X06_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T1_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X06_Y10_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X06_Y10_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X05_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X05_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X06_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X06_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X07_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X07_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X06_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X06_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X06_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X06_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X06_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X06_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T2_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X06_Y10_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X06_Y10_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X05_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X05_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X06_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X06_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X07_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X07_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X06_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X06_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X06_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X06_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X06_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X06_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T3_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X06_Y10_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X06_Y10_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X05_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X05_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X06_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X06_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X07_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X07_Y10_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X06_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X06_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X06_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X06_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X06_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X06_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T4_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X06_Y10_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X06_Y10_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X05_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X05_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X06_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X06_Y10_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y0F_clk_out),
    .clk_out(Tile_X06_Y10_clk_out),
    .clk_pass_through(Tile_X06_Y0F_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X06_Y10_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X06_Y10_clk_pass_through_out_right),
    .config_config_addr(Tile_X06_Y0F_config_out_config_addr),
    .config_config_data(Tile_X06_Y0F_config_out_config_data),
    .config_out_config_addr(Tile_X06_Y10_config_out_config_addr),
    .config_out_config_data(Tile_X06_Y10_config_out_config_data),
    .config_out_read(Tile_X06_Y10_config_out_read),
    .config_out_write(Tile_X06_Y10_config_out_write),
    .config_read(Tile_X06_Y0F_config_out_read),
    .config_write(Tile_X06_Y0F_config_out_write),
    .hi(Tile_X06_Y10_hi),
    .lo(Tile_X06_Y10_lo_unq1),
    .read_config_data(Tile_X06_Y10_read_config_data),
    .read_config_data_in(Tile_X06_Y0F_read_config_data),
    .reset(Tile_X06_Y0F_reset_out),
    .reset_out(Tile_X06_Y10_reset_out),
    .stall(Tile_X06_Y0F_stall_out),
    .stall_out(Tile_X06_Y10_stall_out),
    .tile_id(Tile_X06_Y10_tile_id_in)
);
mantle_wire__typeBit8 Tile_X06_Y10_lo (
    .in(Tile_X06_Y10_lo_unq1),
    .out(Tile_X06_Y10_lo_out)
);
wire [15:0] Tile_X06_Y10_tile_id_out;
assign Tile_X06_Y10_tile_id_out = {Tile_X06_Y10_lo_out[7],Tile_X06_Y10_lo_out[7:6],Tile_X06_Y10_lo_out[6:5],Tile_X06_Y10_hi[5],Tile_X06_Y10_hi[5],Tile_X06_Y10_lo_out[4:3],Tile_X06_Y10_lo_out[3:2],Tile_X06_Y10_hi[2],Tile_X06_Y10_lo_out[1],Tile_X06_Y10_lo_out[1:0],Tile_X06_Y10_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X06_Y10_tile_id (
    .in(Tile_X06_Y10_tile_id_in),
    .out(Tile_X06_Y10_tile_id_out)
);
wire [15:0] Tile_X07_Y00_tile_id;
assign Tile_X07_Y00_tile_id = {Tile_X07_Y00_lo[7],Tile_X07_Y00_lo[7:6],Tile_X07_Y00_lo[6:5],Tile_X07_Y00_hi[5],Tile_X07_Y00_hi[5:4],Tile_X07_Y00_lo[3],Tile_X07_Y00_lo[3:2],Tile_X07_Y00_lo[2:1],Tile_X07_Y00_lo[1:0],Tile_X07_Y00_lo[0]};
Tile_io_core Tile_X07_Y00 (
    .tile_id(Tile_X07_Y00_tile_id),
    .glb2io_1(glb2io_1_X07_Y00),
    .f2io_1(Tile_X07_Y01_SB_T0_NORTH_SB_OUT_B1),
    .io2glb_1(Tile_X07_Y00_io2glb_1),
    .io2f_1(Tile_X07_Y00_io2f_1),
    .glb2io_16(glb2io_16_X07_Y00),
    .f2io_16(Tile_X07_Y01_SB_T0_NORTH_SB_OUT_B16),
    .io2glb_16(Tile_X07_Y00_io2glb_16),
    .io2f_16(Tile_X07_Y00_io2f_16),
    .hi(Tile_X07_Y00_hi),
    .lo(Tile_X07_Y00_lo)
);
Tile_MemCore Tile_X07_Y01 (
    .SB_T0_EAST_SB_IN_B1(Tile_X08_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X08_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X07_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X07_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X07_Y00_io2f_1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X07_Y00_io2f_16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X07_Y01_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X07_Y01_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X07_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X07_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X07_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X07_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X06_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X06_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X07_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X07_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X08_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X08_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X07_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X07_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X07_Y00_io2f_1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X07_Y00_io2f_16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X07_Y01_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X07_Y01_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X07_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X07_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X07_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X07_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X06_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X06_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X07_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X07_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X08_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X08_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X07_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X07_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X07_Y00_io2f_1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X07_Y00_io2f_16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X07_Y01_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X07_Y01_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X07_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X07_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X07_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X07_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X06_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X06_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X07_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X07_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X08_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X08_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X07_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X07_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X07_Y00_io2f_1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X07_Y00_io2f_16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X07_Y01_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X07_Y01_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X07_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X07_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X07_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X07_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X06_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X06_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X07_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X07_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X08_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X08_Y01_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X07_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X07_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X07_Y00_io2f_1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X07_Y00_io2f_16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X07_Y01_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X07_Y01_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X07_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X07_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X07_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X07_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X06_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X06_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X07_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X07_Y01_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y01_clk_pass_through_out_right),
    .clk_out(Tile_X07_Y01_clk_out),
    .config_config_addr(config_7_config_addr),
    .config_config_data(config_7_config_data),
    .config_out_config_addr(Tile_X07_Y01_config_out_config_addr),
    .config_out_config_data(Tile_X07_Y01_config_out_config_data),
    .config_out_read(Tile_X07_Y01_config_out_read),
    .config_out_write(Tile_X07_Y01_config_out_write),
    .config_read(config_7_read),
    .config_write(config_7_write),
    .hi(Tile_X07_Y01_hi_unq1),
    .lo(Tile_X07_Y01_lo_unq1),
    .read_config_data(Tile_X07_Y01_read_config_data),
    .read_config_data_in(const_0_32_out),
    .reset(reset),
    .reset_out(Tile_X07_Y01_reset_out),
    .stall(stall[7]),
    .stall_out(Tile_X07_Y01_stall_out),
    .tile_id(Tile_X07_Y01_tile_id_in)
);
mantle_wire__typeBit9 Tile_X07_Y01_hi (
    .in(Tile_X07_Y01_hi_unq1),
    .out(Tile_X07_Y01_hi_out)
);
mantle_wire__typeBit8 Tile_X07_Y01_lo (
    .in(Tile_X07_Y01_lo_unq1),
    .out(Tile_X07_Y01_lo_out)
);
wire [15:0] Tile_X07_Y01_tile_id_out;
assign Tile_X07_Y01_tile_id_out = {Tile_X07_Y01_lo_out[7],Tile_X07_Y01_lo_out[7:6],Tile_X07_Y01_lo_out[6:5],Tile_X07_Y01_hi_out[5],Tile_X07_Y01_hi_out[5:4],Tile_X07_Y01_lo_out[3],Tile_X07_Y01_lo_out[3:2],Tile_X07_Y01_lo_out[2:1],Tile_X07_Y01_lo_out[1:0],Tile_X07_Y01_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X07_Y01_tile_id (
    .in(Tile_X07_Y01_tile_id_in),
    .out(Tile_X07_Y01_tile_id_out)
);
Tile_MemCore Tile_X07_Y02 (
    .SB_T0_EAST_SB_IN_B1(Tile_X08_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X08_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X07_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X07_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X07_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X07_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X07_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X07_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X07_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X07_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X07_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X07_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X06_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X06_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X07_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X07_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X08_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X08_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X07_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X07_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X07_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X07_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X07_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X07_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X07_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X07_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X07_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X07_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X06_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X06_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X07_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X07_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X08_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X08_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X07_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X07_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X07_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X07_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X07_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X07_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X07_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X07_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X07_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X07_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X06_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X06_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X07_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X07_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X08_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X08_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X07_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X07_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X07_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X07_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X07_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X07_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X07_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X07_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X07_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X07_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X06_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X06_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X07_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X07_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X08_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X08_Y02_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X07_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X07_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X07_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X07_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X07_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X07_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X07_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X07_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X07_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X07_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X06_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X06_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X07_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X07_Y02_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y02_clk_pass_through_out_right),
    .clk_out(Tile_X07_Y02_clk_out),
    .config_config_addr(Tile_X07_Y01_config_out_config_addr),
    .config_config_data(Tile_X07_Y01_config_out_config_data),
    .config_out_config_addr(Tile_X07_Y02_config_out_config_addr),
    .config_out_config_data(Tile_X07_Y02_config_out_config_data),
    .config_out_read(Tile_X07_Y02_config_out_read),
    .config_out_write(Tile_X07_Y02_config_out_write),
    .config_read(Tile_X07_Y01_config_out_read),
    .config_write(Tile_X07_Y01_config_out_write),
    .hi(Tile_X07_Y02_hi_unq1),
    .lo(Tile_X07_Y02_lo_unq1),
    .read_config_data(Tile_X07_Y02_read_config_data),
    .read_config_data_in(Tile_X07_Y01_read_config_data),
    .reset(Tile_X07_Y01_reset_out),
    .reset_out(Tile_X07_Y02_reset_out),
    .stall(Tile_X07_Y01_stall_out),
    .stall_out(Tile_X07_Y02_stall_out),
    .tile_id(Tile_X07_Y02_tile_id_in)
);
mantle_wire__typeBit9 Tile_X07_Y02_hi (
    .in(Tile_X07_Y02_hi_unq1),
    .out(Tile_X07_Y02_hi_out)
);
mantle_wire__typeBit8 Tile_X07_Y02_lo (
    .in(Tile_X07_Y02_lo_unq1),
    .out(Tile_X07_Y02_lo_out)
);
wire [15:0] Tile_X07_Y02_tile_id_out;
assign Tile_X07_Y02_tile_id_out = {Tile_X07_Y02_lo_out[7],Tile_X07_Y02_lo_out[7:6],Tile_X07_Y02_lo_out[6:5],Tile_X07_Y02_hi_out[5],Tile_X07_Y02_hi_out[5:4],Tile_X07_Y02_lo_out[3],Tile_X07_Y02_lo_out[3:2],Tile_X07_Y02_lo_out[2:1],Tile_X07_Y02_lo_out[1],Tile_X07_Y02_hi_out[1],Tile_X07_Y02_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X07_Y02_tile_id (
    .in(Tile_X07_Y02_tile_id_in),
    .out(Tile_X07_Y02_tile_id_out)
);
Tile_MemCore Tile_X07_Y03 (
    .SB_T0_EAST_SB_IN_B1(Tile_X08_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X08_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X07_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X07_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X07_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X07_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X07_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X07_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X07_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X07_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X07_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X07_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X06_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X06_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X07_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X07_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X08_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X08_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X07_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X07_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X07_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X07_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X07_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X07_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X07_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X07_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X07_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X07_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X06_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X06_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X07_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X07_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X08_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X08_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X07_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X07_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X07_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X07_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X07_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X07_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X07_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X07_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X07_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X07_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X06_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X06_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X07_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X07_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X08_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X08_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X07_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X07_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X07_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X07_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X07_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X07_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X07_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X07_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X07_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X07_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X06_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X06_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X07_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X07_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X08_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X08_Y03_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X07_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X07_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X07_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X07_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X07_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X07_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X07_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X07_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X07_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X07_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X06_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X06_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X07_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X07_Y03_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y03_clk_pass_through_out_right),
    .clk_out(Tile_X07_Y03_clk_out),
    .config_config_addr(Tile_X07_Y02_config_out_config_addr),
    .config_config_data(Tile_X07_Y02_config_out_config_data),
    .config_out_config_addr(Tile_X07_Y03_config_out_config_addr),
    .config_out_config_data(Tile_X07_Y03_config_out_config_data),
    .config_out_read(Tile_X07_Y03_config_out_read),
    .config_out_write(Tile_X07_Y03_config_out_write),
    .config_read(Tile_X07_Y02_config_out_read),
    .config_write(Tile_X07_Y02_config_out_write),
    .hi(Tile_X07_Y03_hi_unq1),
    .lo(Tile_X07_Y03_lo_unq1),
    .read_config_data(Tile_X07_Y03_read_config_data),
    .read_config_data_in(Tile_X07_Y02_read_config_data),
    .reset(Tile_X07_Y02_reset_out),
    .reset_out(Tile_X07_Y03_reset_out),
    .stall(Tile_X07_Y02_stall_out),
    .stall_out(Tile_X07_Y03_stall_out),
    .tile_id(Tile_X07_Y03_tile_id_in)
);
mantle_wire__typeBit9 Tile_X07_Y03_hi (
    .in(Tile_X07_Y03_hi_unq1),
    .out(Tile_X07_Y03_hi_out)
);
mantle_wire__typeBit8 Tile_X07_Y03_lo (
    .in(Tile_X07_Y03_lo_unq1),
    .out(Tile_X07_Y03_lo_out)
);
wire [15:0] Tile_X07_Y03_tile_id_out;
assign Tile_X07_Y03_tile_id_out = {Tile_X07_Y03_lo_out[7],Tile_X07_Y03_lo_out[7:6],Tile_X07_Y03_lo_out[6:5],Tile_X07_Y03_hi_out[5],Tile_X07_Y03_hi_out[5:4],Tile_X07_Y03_lo_out[3],Tile_X07_Y03_lo_out[3:2],Tile_X07_Y03_lo_out[2:1],Tile_X07_Y03_lo_out[1],Tile_X07_Y03_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X07_Y03_tile_id (
    .in(Tile_X07_Y03_tile_id_in),
    .out(Tile_X07_Y03_tile_id_out)
);
Tile_MemCore Tile_X07_Y04 (
    .SB_T0_EAST_SB_IN_B1(Tile_X08_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X08_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X07_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X07_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X07_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X07_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X07_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X07_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X07_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X07_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X07_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X07_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X06_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X06_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X07_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X07_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X08_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X08_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X07_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X07_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X07_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X07_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X07_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X07_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X07_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X07_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X07_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X07_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X06_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X06_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X07_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X07_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X08_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X08_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X07_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X07_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X07_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X07_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X07_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X07_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X07_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X07_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X07_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X07_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X06_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X06_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X07_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X07_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X08_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X08_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X07_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X07_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X07_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X07_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X07_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X07_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X07_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X07_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X07_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X07_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X06_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X06_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X07_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X07_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X08_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X08_Y04_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X07_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X07_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X07_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X07_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X07_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X07_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X07_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X07_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X07_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X07_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X06_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X06_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X07_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X07_Y04_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y04_clk_pass_through_out_right),
    .clk_out(Tile_X07_Y04_clk_out),
    .config_config_addr(Tile_X07_Y03_config_out_config_addr),
    .config_config_data(Tile_X07_Y03_config_out_config_data),
    .config_out_config_addr(Tile_X07_Y04_config_out_config_addr),
    .config_out_config_data(Tile_X07_Y04_config_out_config_data),
    .config_out_read(Tile_X07_Y04_config_out_read),
    .config_out_write(Tile_X07_Y04_config_out_write),
    .config_read(Tile_X07_Y03_config_out_read),
    .config_write(Tile_X07_Y03_config_out_write),
    .hi(Tile_X07_Y04_hi_unq1),
    .lo(Tile_X07_Y04_lo_unq1),
    .read_config_data(Tile_X07_Y04_read_config_data),
    .read_config_data_in(Tile_X07_Y03_read_config_data),
    .reset(Tile_X07_Y03_reset_out),
    .reset_out(Tile_X07_Y04_reset_out),
    .stall(Tile_X07_Y03_stall_out),
    .stall_out(Tile_X07_Y04_stall_out),
    .tile_id(Tile_X07_Y04_tile_id_in)
);
mantle_wire__typeBit9 Tile_X07_Y04_hi (
    .in(Tile_X07_Y04_hi_unq1),
    .out(Tile_X07_Y04_hi_out)
);
mantle_wire__typeBit8 Tile_X07_Y04_lo (
    .in(Tile_X07_Y04_lo_unq1),
    .out(Tile_X07_Y04_lo_out)
);
wire [15:0] Tile_X07_Y04_tile_id_out;
assign Tile_X07_Y04_tile_id_out = {Tile_X07_Y04_lo_out[7],Tile_X07_Y04_lo_out[7:6],Tile_X07_Y04_lo_out[6:5],Tile_X07_Y04_hi_out[5],Tile_X07_Y04_hi_out[5:4],Tile_X07_Y04_lo_out[3],Tile_X07_Y04_lo_out[3:2],Tile_X07_Y04_lo_out[2:1],Tile_X07_Y04_hi_out[1],Tile_X07_Y04_lo_out[0],Tile_X07_Y04_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X07_Y04_tile_id (
    .in(Tile_X07_Y04_tile_id_in),
    .out(Tile_X07_Y04_tile_id_out)
);
Tile_MemCore Tile_X07_Y05 (
    .SB_T0_EAST_SB_IN_B1(Tile_X08_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X08_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X07_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X07_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X07_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X07_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X07_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X07_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X07_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X07_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X07_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X07_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X06_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X06_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X07_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X07_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X08_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X08_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X07_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X07_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X07_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X07_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X07_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X07_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X07_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X07_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X07_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X07_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X06_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X06_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X07_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X07_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X08_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X08_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X07_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X07_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X07_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X07_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X07_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X07_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X07_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X07_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X07_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X07_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X06_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X06_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X07_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X07_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X08_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X08_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X07_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X07_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X07_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X07_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X07_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X07_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X07_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X07_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X07_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X07_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X06_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X06_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X07_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X07_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X08_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X08_Y05_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X07_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X07_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X07_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X07_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X07_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X07_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X07_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X07_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X07_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X07_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X06_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X06_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X07_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X07_Y05_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y05_clk_pass_through_out_right),
    .clk_out(Tile_X07_Y05_clk_out),
    .config_config_addr(Tile_X07_Y04_config_out_config_addr),
    .config_config_data(Tile_X07_Y04_config_out_config_data),
    .config_out_config_addr(Tile_X07_Y05_config_out_config_addr),
    .config_out_config_data(Tile_X07_Y05_config_out_config_data),
    .config_out_read(Tile_X07_Y05_config_out_read),
    .config_out_write(Tile_X07_Y05_config_out_write),
    .config_read(Tile_X07_Y04_config_out_read),
    .config_write(Tile_X07_Y04_config_out_write),
    .hi(Tile_X07_Y05_hi_unq1),
    .lo(Tile_X07_Y05_lo_unq1),
    .read_config_data(Tile_X07_Y05_read_config_data),
    .read_config_data_in(Tile_X07_Y04_read_config_data),
    .reset(Tile_X07_Y04_reset_out),
    .reset_out(Tile_X07_Y05_reset_out),
    .stall(Tile_X07_Y04_stall_out),
    .stall_out(Tile_X07_Y05_stall_out),
    .tile_id(Tile_X07_Y05_tile_id_in)
);
mantle_wire__typeBit9 Tile_X07_Y05_hi (
    .in(Tile_X07_Y05_hi_unq1),
    .out(Tile_X07_Y05_hi_out)
);
mantle_wire__typeBit8 Tile_X07_Y05_lo (
    .in(Tile_X07_Y05_lo_unq1),
    .out(Tile_X07_Y05_lo_out)
);
wire [15:0] Tile_X07_Y05_tile_id_out;
assign Tile_X07_Y05_tile_id_out = {Tile_X07_Y05_lo_out[7],Tile_X07_Y05_lo_out[7:6],Tile_X07_Y05_lo_out[6:5],Tile_X07_Y05_hi_out[5],Tile_X07_Y05_hi_out[5:4],Tile_X07_Y05_lo_out[3],Tile_X07_Y05_lo_out[3:2],Tile_X07_Y05_lo_out[2:1],Tile_X07_Y05_hi_out[1],Tile_X07_Y05_lo_out[0],Tile_X07_Y05_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X07_Y05_tile_id (
    .in(Tile_X07_Y05_tile_id_in),
    .out(Tile_X07_Y05_tile_id_out)
);
Tile_MemCore Tile_X07_Y06 (
    .SB_T0_EAST_SB_IN_B1(Tile_X08_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X08_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X07_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X07_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X07_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X07_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X07_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X07_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X07_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X07_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X07_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X07_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X06_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X06_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X07_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X07_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X08_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X08_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X07_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X07_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X07_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X07_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X07_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X07_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X07_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X07_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X07_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X07_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X06_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X06_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X07_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X07_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X08_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X08_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X07_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X07_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X07_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X07_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X07_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X07_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X07_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X07_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X07_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X07_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X06_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X06_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X07_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X07_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X08_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X08_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X07_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X07_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X07_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X07_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X07_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X07_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X07_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X07_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X07_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X07_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X06_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X06_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X07_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X07_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X08_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X08_Y06_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X07_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X07_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X07_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X07_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X07_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X07_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X07_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X07_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X07_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X07_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X06_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X06_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X07_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X07_Y06_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y06_clk_pass_through_out_right),
    .clk_out(Tile_X07_Y06_clk_out),
    .config_config_addr(Tile_X07_Y05_config_out_config_addr),
    .config_config_data(Tile_X07_Y05_config_out_config_data),
    .config_out_config_addr(Tile_X07_Y06_config_out_config_addr),
    .config_out_config_data(Tile_X07_Y06_config_out_config_data),
    .config_out_read(Tile_X07_Y06_config_out_read),
    .config_out_write(Tile_X07_Y06_config_out_write),
    .config_read(Tile_X07_Y05_config_out_read),
    .config_write(Tile_X07_Y05_config_out_write),
    .hi(Tile_X07_Y06_hi_unq1),
    .lo(Tile_X07_Y06_lo_unq1),
    .read_config_data(Tile_X07_Y06_read_config_data),
    .read_config_data_in(Tile_X07_Y05_read_config_data),
    .reset(Tile_X07_Y05_reset_out),
    .reset_out(Tile_X07_Y06_reset_out),
    .stall(Tile_X07_Y05_stall_out),
    .stall_out(Tile_X07_Y06_stall_out),
    .tile_id(Tile_X07_Y06_tile_id_in)
);
mantle_wire__typeBit9 Tile_X07_Y06_hi (
    .in(Tile_X07_Y06_hi_unq1),
    .out(Tile_X07_Y06_hi_out)
);
mantle_wire__typeBit8 Tile_X07_Y06_lo (
    .in(Tile_X07_Y06_lo_unq1),
    .out(Tile_X07_Y06_lo_out)
);
wire [15:0] Tile_X07_Y06_tile_id_out;
assign Tile_X07_Y06_tile_id_out = {Tile_X07_Y06_lo_out[7],Tile_X07_Y06_lo_out[7:6],Tile_X07_Y06_lo_out[6:5],Tile_X07_Y06_hi_out[5],Tile_X07_Y06_hi_out[5:4],Tile_X07_Y06_lo_out[3],Tile_X07_Y06_lo_out[3:2],Tile_X07_Y06_lo_out[2:1],Tile_X07_Y06_hi_out[1],Tile_X07_Y06_hi_out[1],Tile_X07_Y06_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X07_Y06_tile_id (
    .in(Tile_X07_Y06_tile_id_in),
    .out(Tile_X07_Y06_tile_id_out)
);
Tile_MemCore Tile_X07_Y07 (
    .SB_T0_EAST_SB_IN_B1(Tile_X08_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X08_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X07_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X07_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X07_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X07_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X07_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X07_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X07_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X07_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X07_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X07_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X06_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X06_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X07_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X07_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X08_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X08_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X07_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X07_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X07_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X07_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X07_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X07_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X07_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X07_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X07_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X07_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X06_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X06_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X07_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X07_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X08_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X08_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X07_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X07_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X07_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X07_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X07_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X07_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X07_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X07_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X07_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X07_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X06_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X06_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X07_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X07_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X08_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X08_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X07_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X07_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X07_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X07_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X07_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X07_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X07_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X07_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X07_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X07_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X06_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X06_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X07_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X07_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X08_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X08_Y07_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X07_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X07_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X07_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X07_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X07_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X07_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X07_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X07_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X07_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X07_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X06_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X06_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X07_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X07_Y07_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y07_clk_pass_through_out_right),
    .clk_out(Tile_X07_Y07_clk_out),
    .config_config_addr(Tile_X07_Y06_config_out_config_addr),
    .config_config_data(Tile_X07_Y06_config_out_config_data),
    .config_out_config_addr(Tile_X07_Y07_config_out_config_addr),
    .config_out_config_data(Tile_X07_Y07_config_out_config_data),
    .config_out_read(Tile_X07_Y07_config_out_read),
    .config_out_write(Tile_X07_Y07_config_out_write),
    .config_read(Tile_X07_Y06_config_out_read),
    .config_write(Tile_X07_Y06_config_out_write),
    .hi(Tile_X07_Y07_hi_unq1),
    .lo(Tile_X07_Y07_lo_unq1),
    .read_config_data(Tile_X07_Y07_read_config_data),
    .read_config_data_in(Tile_X07_Y06_read_config_data),
    .reset(Tile_X07_Y06_reset_out),
    .reset_out(Tile_X07_Y07_reset_out),
    .stall(Tile_X07_Y06_stall_out),
    .stall_out(Tile_X07_Y07_stall_out),
    .tile_id(Tile_X07_Y07_tile_id_in)
);
mantle_wire__typeBit9 Tile_X07_Y07_hi (
    .in(Tile_X07_Y07_hi_unq1),
    .out(Tile_X07_Y07_hi_out)
);
mantle_wire__typeBit8 Tile_X07_Y07_lo (
    .in(Tile_X07_Y07_lo_unq1),
    .out(Tile_X07_Y07_lo_out)
);
wire [15:0] Tile_X07_Y07_tile_id_out;
assign Tile_X07_Y07_tile_id_out = {Tile_X07_Y07_lo_out[7],Tile_X07_Y07_lo_out[7:6],Tile_X07_Y07_lo_out[6:5],Tile_X07_Y07_hi_out[5],Tile_X07_Y07_hi_out[5:4],Tile_X07_Y07_lo_out[3],Tile_X07_Y07_lo_out[3:2],Tile_X07_Y07_lo_out[2:1],Tile_X07_Y07_hi_out[1],Tile_X07_Y07_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X07_Y07_tile_id (
    .in(Tile_X07_Y07_tile_id_in),
    .out(Tile_X07_Y07_tile_id_out)
);
Tile_MemCore Tile_X07_Y08 (
    .SB_T0_EAST_SB_IN_B1(Tile_X08_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X08_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X07_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X07_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X07_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X07_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X07_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X07_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X07_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X07_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X07_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X07_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X06_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X06_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X07_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X07_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X08_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X08_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X07_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X07_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X07_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X07_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X07_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X07_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X07_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X07_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X07_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X07_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X06_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X06_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X07_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X07_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X08_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X08_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X07_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X07_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X07_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X07_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X07_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X07_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X07_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X07_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X07_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X07_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X06_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X06_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X07_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X07_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X08_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X08_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X07_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X07_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X07_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X07_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X07_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X07_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X07_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X07_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X07_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X07_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X06_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X06_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X07_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X07_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X08_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X08_Y08_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X07_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X07_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X07_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X07_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X07_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X07_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X07_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X07_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X07_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X07_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X06_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X06_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X07_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X07_Y08_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y08_clk_pass_through_out_right),
    .clk_out(Tile_X07_Y08_clk_out),
    .config_config_addr(Tile_X07_Y07_config_out_config_addr),
    .config_config_data(Tile_X07_Y07_config_out_config_data),
    .config_out_config_addr(Tile_X07_Y08_config_out_config_addr),
    .config_out_config_data(Tile_X07_Y08_config_out_config_data),
    .config_out_read(Tile_X07_Y08_config_out_read),
    .config_out_write(Tile_X07_Y08_config_out_write),
    .config_read(Tile_X07_Y07_config_out_read),
    .config_write(Tile_X07_Y07_config_out_write),
    .hi(Tile_X07_Y08_hi_unq1),
    .lo(Tile_X07_Y08_lo_unq1),
    .read_config_data(Tile_X07_Y08_read_config_data),
    .read_config_data_in(Tile_X07_Y07_read_config_data),
    .reset(Tile_X07_Y07_reset_out),
    .reset_out(Tile_X07_Y08_reset_out),
    .stall(Tile_X07_Y07_stall_out),
    .stall_out(Tile_X07_Y08_stall_out),
    .tile_id(Tile_X07_Y08_tile_id_in)
);
mantle_wire__typeBit9 Tile_X07_Y08_hi (
    .in(Tile_X07_Y08_hi_unq1),
    .out(Tile_X07_Y08_hi_out)
);
mantle_wire__typeBit8 Tile_X07_Y08_lo (
    .in(Tile_X07_Y08_lo_unq1),
    .out(Tile_X07_Y08_lo_out)
);
wire [15:0] Tile_X07_Y08_tile_id_out;
assign Tile_X07_Y08_tile_id_out = {Tile_X07_Y08_lo_out[7],Tile_X07_Y08_lo_out[7:6],Tile_X07_Y08_lo_out[6:5],Tile_X07_Y08_hi_out[5],Tile_X07_Y08_hi_out[5:4],Tile_X07_Y08_lo_out[3],Tile_X07_Y08_lo_out[3:2],Tile_X07_Y08_lo_out[2],Tile_X07_Y08_hi_out[2],Tile_X07_Y08_lo_out[1:0],Tile_X07_Y08_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X07_Y08_tile_id (
    .in(Tile_X07_Y08_tile_id_in),
    .out(Tile_X07_Y08_tile_id_out)
);
Tile_MemCore Tile_X07_Y09 (
    .SB_T0_EAST_SB_IN_B1(Tile_X08_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X08_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X07_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X07_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X07_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X07_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X07_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X07_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X07_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X07_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X07_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X07_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X06_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X06_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X07_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X07_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X08_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X08_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X07_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X07_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X07_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X07_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X07_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X07_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X07_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X07_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X07_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X07_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X06_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X06_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X07_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X07_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X08_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X08_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X07_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X07_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X07_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X07_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X07_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X07_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X07_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X07_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X07_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X07_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X06_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X06_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X07_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X07_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X08_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X08_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X07_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X07_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X07_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X07_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X07_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X07_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X07_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X07_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X07_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X07_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X06_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X06_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X07_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X07_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X08_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X08_Y09_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X07_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X07_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X07_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X07_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X07_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X07_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X07_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X07_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X07_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X07_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X06_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X06_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X07_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X07_Y09_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y09_clk_pass_through_out_right),
    .clk_out(Tile_X07_Y09_clk_out),
    .config_config_addr(ConfigPipeStage_inst7_config_out_config_addr),
    .config_config_data(ConfigPipeStage_inst7_config_out_config_data),
    .config_out_config_addr(Tile_X07_Y09_config_out_config_addr),
    .config_out_config_data(Tile_X07_Y09_config_out_config_data),
    .config_out_read(Tile_X07_Y09_config_out_read),
    .config_out_write(Tile_X07_Y09_config_out_write),
    .config_read(ConfigPipeStage_inst7_config_out_read),
    .config_write(ConfigPipeStage_inst7_config_out_write),
    .hi(Tile_X07_Y09_hi_unq1),
    .lo(Tile_X07_Y09_lo_unq1),
    .read_config_data(Tile_X07_Y09_read_config_data),
    .read_config_data_in(Tile_X07_Y08_read_config_data),
    .reset(Tile_X07_Y08_reset_out),
    .reset_out(Tile_X07_Y09_reset_out),
    .stall(Tile_X07_Y08_stall_out),
    .stall_out(Tile_X07_Y09_stall_out),
    .tile_id(Tile_X07_Y09_tile_id_in)
);
mantle_wire__typeBit9 Tile_X07_Y09_hi (
    .in(Tile_X07_Y09_hi_unq1),
    .out(Tile_X07_Y09_hi_out)
);
mantle_wire__typeBit8 Tile_X07_Y09_lo (
    .in(Tile_X07_Y09_lo_unq1),
    .out(Tile_X07_Y09_lo_out)
);
wire [15:0] Tile_X07_Y09_tile_id_out;
assign Tile_X07_Y09_tile_id_out = {Tile_X07_Y09_lo_out[7],Tile_X07_Y09_lo_out[7:6],Tile_X07_Y09_lo_out[6:5],Tile_X07_Y09_hi_out[5],Tile_X07_Y09_hi_out[5:4],Tile_X07_Y09_lo_out[3],Tile_X07_Y09_lo_out[3:2],Tile_X07_Y09_lo_out[2],Tile_X07_Y09_hi_out[2],Tile_X07_Y09_lo_out[1:0],Tile_X07_Y09_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X07_Y09_tile_id (
    .in(Tile_X07_Y09_tile_id_in),
    .out(Tile_X07_Y09_tile_id_out)
);
Tile_MemCore Tile_X07_Y0A (
    .SB_T0_EAST_SB_IN_B1(Tile_X08_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X08_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X07_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X07_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X07_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X07_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X07_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X07_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X07_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X07_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X07_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X07_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X06_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X06_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X07_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X07_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X08_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X08_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X07_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X07_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X07_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X07_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X07_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X07_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X07_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X07_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X07_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X07_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X06_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X06_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X07_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X07_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X08_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X08_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X07_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X07_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X07_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X07_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X07_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X07_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X07_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X07_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X07_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X07_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X06_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X06_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X07_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X07_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X08_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X08_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X07_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X07_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X07_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X07_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X07_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X07_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X07_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X07_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X07_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X07_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X06_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X06_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X07_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X07_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X08_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X08_Y0A_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X07_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X07_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X07_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X07_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X07_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X07_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X07_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X07_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X07_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X07_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X06_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X06_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X07_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X07_Y0A_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y0A_clk_pass_through_out_right),
    .clk_out(Tile_X07_Y0A_clk_out),
    .config_config_addr(Tile_X07_Y09_config_out_config_addr),
    .config_config_data(Tile_X07_Y09_config_out_config_data),
    .config_out_config_addr(Tile_X07_Y0A_config_out_config_addr),
    .config_out_config_data(Tile_X07_Y0A_config_out_config_data),
    .config_out_read(Tile_X07_Y0A_config_out_read),
    .config_out_write(Tile_X07_Y0A_config_out_write),
    .config_read(Tile_X07_Y09_config_out_read),
    .config_write(Tile_X07_Y09_config_out_write),
    .hi(Tile_X07_Y0A_hi_unq1),
    .lo(Tile_X07_Y0A_lo_unq1),
    .read_config_data(Tile_X07_Y0A_read_config_data),
    .read_config_data_in(Tile_X07_Y09_read_config_data),
    .reset(Tile_X07_Y09_reset_out),
    .reset_out(Tile_X07_Y0A_reset_out),
    .stall(Tile_X07_Y09_stall_out),
    .stall_out(Tile_X07_Y0A_stall_out),
    .tile_id(Tile_X07_Y0A_tile_id_in)
);
mantle_wire__typeBit9 Tile_X07_Y0A_hi (
    .in(Tile_X07_Y0A_hi_unq1),
    .out(Tile_X07_Y0A_hi_out)
);
mantle_wire__typeBit8 Tile_X07_Y0A_lo (
    .in(Tile_X07_Y0A_lo_unq1),
    .out(Tile_X07_Y0A_lo_out)
);
wire [15:0] Tile_X07_Y0A_tile_id_out;
assign Tile_X07_Y0A_tile_id_out = {Tile_X07_Y0A_lo_out[7],Tile_X07_Y0A_lo_out[7:6],Tile_X07_Y0A_lo_out[6:5],Tile_X07_Y0A_hi_out[5],Tile_X07_Y0A_hi_out[5:4],Tile_X07_Y0A_lo_out[3],Tile_X07_Y0A_lo_out[3:2],Tile_X07_Y0A_lo_out[2],Tile_X07_Y0A_hi_out[2],Tile_X07_Y0A_lo_out[1],Tile_X07_Y0A_hi_out[1],Tile_X07_Y0A_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X07_Y0A_tile_id (
    .in(Tile_X07_Y0A_tile_id_in),
    .out(Tile_X07_Y0A_tile_id_out)
);
Tile_MemCore Tile_X07_Y0B (
    .SB_T0_EAST_SB_IN_B1(Tile_X08_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X08_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X07_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X07_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X07_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X07_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X07_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X07_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X07_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X07_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X07_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X07_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X06_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X06_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X07_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X07_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X08_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X08_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X07_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X07_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X07_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X07_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X07_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X07_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X07_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X07_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X07_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X07_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X06_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X06_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X07_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X07_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X08_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X08_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X07_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X07_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X07_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X07_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X07_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X07_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X07_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X07_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X07_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X07_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X06_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X06_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X07_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X07_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X08_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X08_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X07_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X07_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X07_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X07_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X07_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X07_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X07_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X07_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X07_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X07_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X06_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X06_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X07_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X07_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X08_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X08_Y0B_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X07_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X07_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X07_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X07_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X07_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X07_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X07_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X07_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X07_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X07_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X06_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X06_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X07_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X07_Y0B_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y0B_clk_pass_through_out_right),
    .clk_out(Tile_X07_Y0B_clk_out),
    .config_config_addr(Tile_X07_Y0A_config_out_config_addr),
    .config_config_data(Tile_X07_Y0A_config_out_config_data),
    .config_out_config_addr(Tile_X07_Y0B_config_out_config_addr),
    .config_out_config_data(Tile_X07_Y0B_config_out_config_data),
    .config_out_read(Tile_X07_Y0B_config_out_read),
    .config_out_write(Tile_X07_Y0B_config_out_write),
    .config_read(Tile_X07_Y0A_config_out_read),
    .config_write(Tile_X07_Y0A_config_out_write),
    .hi(Tile_X07_Y0B_hi_unq1),
    .lo(Tile_X07_Y0B_lo_unq1),
    .read_config_data(Tile_X07_Y0B_read_config_data),
    .read_config_data_in(Tile_X07_Y0A_read_config_data),
    .reset(Tile_X07_Y0A_reset_out),
    .reset_out(Tile_X07_Y0B_reset_out),
    .stall(Tile_X07_Y0A_stall_out),
    .stall_out(Tile_X07_Y0B_stall_out),
    .tile_id(Tile_X07_Y0B_tile_id_in)
);
mantle_wire__typeBit9 Tile_X07_Y0B_hi (
    .in(Tile_X07_Y0B_hi_unq1),
    .out(Tile_X07_Y0B_hi_out)
);
mantle_wire__typeBit8 Tile_X07_Y0B_lo (
    .in(Tile_X07_Y0B_lo_unq1),
    .out(Tile_X07_Y0B_lo_out)
);
wire [15:0] Tile_X07_Y0B_tile_id_out;
assign Tile_X07_Y0B_tile_id_out = {Tile_X07_Y0B_lo_out[7],Tile_X07_Y0B_lo_out[7:6],Tile_X07_Y0B_lo_out[6:5],Tile_X07_Y0B_hi_out[5],Tile_X07_Y0B_hi_out[5:4],Tile_X07_Y0B_lo_out[3],Tile_X07_Y0B_lo_out[3:2],Tile_X07_Y0B_lo_out[2],Tile_X07_Y0B_hi_out[2],Tile_X07_Y0B_lo_out[1],Tile_X07_Y0B_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X07_Y0B_tile_id (
    .in(Tile_X07_Y0B_tile_id_in),
    .out(Tile_X07_Y0B_tile_id_out)
);
Tile_MemCore Tile_X07_Y0C (
    .SB_T0_EAST_SB_IN_B1(Tile_X08_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X08_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X07_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X07_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X07_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X07_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X07_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X07_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X07_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X07_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X07_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X07_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X06_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X06_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X07_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X07_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X08_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X08_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X07_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X07_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X07_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X07_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X07_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X07_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X07_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X07_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X07_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X07_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X06_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X06_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X07_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X07_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X08_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X08_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X07_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X07_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X07_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X07_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X07_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X07_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X07_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X07_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X07_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X07_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X06_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X06_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X07_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X07_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X08_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X08_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X07_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X07_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X07_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X07_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X07_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X07_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X07_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X07_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X07_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X07_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X06_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X06_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X07_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X07_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X08_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X08_Y0C_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X07_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X07_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X07_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X07_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X07_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X07_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X07_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X07_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X07_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X07_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X06_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X06_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X07_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X07_Y0C_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y0C_clk_pass_through_out_right),
    .clk_out(Tile_X07_Y0C_clk_out),
    .config_config_addr(Tile_X07_Y0B_config_out_config_addr),
    .config_config_data(Tile_X07_Y0B_config_out_config_data),
    .config_out_config_addr(Tile_X07_Y0C_config_out_config_addr),
    .config_out_config_data(Tile_X07_Y0C_config_out_config_data),
    .config_out_read(Tile_X07_Y0C_config_out_read),
    .config_out_write(Tile_X07_Y0C_config_out_write),
    .config_read(Tile_X07_Y0B_config_out_read),
    .config_write(Tile_X07_Y0B_config_out_write),
    .hi(Tile_X07_Y0C_hi_unq1),
    .lo(Tile_X07_Y0C_lo_unq1),
    .read_config_data(Tile_X07_Y0C_read_config_data),
    .read_config_data_in(Tile_X07_Y0B_read_config_data),
    .reset(Tile_X07_Y0B_reset_out),
    .reset_out(Tile_X07_Y0C_reset_out),
    .stall(Tile_X07_Y0B_stall_out),
    .stall_out(Tile_X07_Y0C_stall_out),
    .tile_id(Tile_X07_Y0C_tile_id_in)
);
mantle_wire__typeBit9 Tile_X07_Y0C_hi (
    .in(Tile_X07_Y0C_hi_unq1),
    .out(Tile_X07_Y0C_hi_out)
);
mantle_wire__typeBit8 Tile_X07_Y0C_lo (
    .in(Tile_X07_Y0C_lo_unq1),
    .out(Tile_X07_Y0C_lo_out)
);
wire [15:0] Tile_X07_Y0C_tile_id_out;
assign Tile_X07_Y0C_tile_id_out = {Tile_X07_Y0C_lo_out[7],Tile_X07_Y0C_lo_out[7:6],Tile_X07_Y0C_lo_out[6:5],Tile_X07_Y0C_hi_out[5],Tile_X07_Y0C_hi_out[5:4],Tile_X07_Y0C_lo_out[3],Tile_X07_Y0C_lo_out[3:2],Tile_X07_Y0C_lo_out[2],Tile_X07_Y0C_hi_out[2:1],Tile_X07_Y0C_lo_out[0],Tile_X07_Y0C_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X07_Y0C_tile_id (
    .in(Tile_X07_Y0C_tile_id_in),
    .out(Tile_X07_Y0C_tile_id_out)
);
Tile_MemCore Tile_X07_Y0D (
    .SB_T0_EAST_SB_IN_B1(Tile_X08_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X08_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X07_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X07_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X07_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X07_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X07_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X07_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X07_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X07_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X07_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X07_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X06_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X06_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X07_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X07_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X08_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X08_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X07_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X07_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X07_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X07_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X07_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X07_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X07_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X07_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X07_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X07_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X06_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X06_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X07_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X07_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X08_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X08_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X07_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X07_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X07_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X07_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X07_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X07_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X07_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X07_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X07_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X07_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X06_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X06_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X07_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X07_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X08_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X08_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X07_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X07_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X07_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X07_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X07_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X07_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X07_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X07_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X07_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X07_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X06_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X06_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X07_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X07_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X08_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X08_Y0D_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X07_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X07_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X07_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X07_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X07_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X07_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X07_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X07_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X07_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X07_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X06_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X06_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X07_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X07_Y0D_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y0D_clk_pass_through_out_right),
    .clk_out(Tile_X07_Y0D_clk_out),
    .config_config_addr(Tile_X07_Y0C_config_out_config_addr),
    .config_config_data(Tile_X07_Y0C_config_out_config_data),
    .config_out_config_addr(Tile_X07_Y0D_config_out_config_addr),
    .config_out_config_data(Tile_X07_Y0D_config_out_config_data),
    .config_out_read(Tile_X07_Y0D_config_out_read),
    .config_out_write(Tile_X07_Y0D_config_out_write),
    .config_read(Tile_X07_Y0C_config_out_read),
    .config_write(Tile_X07_Y0C_config_out_write),
    .hi(Tile_X07_Y0D_hi_unq1),
    .lo(Tile_X07_Y0D_lo_unq1),
    .read_config_data(Tile_X07_Y0D_read_config_data),
    .read_config_data_in(Tile_X07_Y0C_read_config_data),
    .reset(Tile_X07_Y0C_reset_out),
    .reset_out(Tile_X07_Y0D_reset_out),
    .stall(Tile_X07_Y0C_stall_out),
    .stall_out(Tile_X07_Y0D_stall_out),
    .tile_id(Tile_X07_Y0D_tile_id_in)
);
mantle_wire__typeBit9 Tile_X07_Y0D_hi (
    .in(Tile_X07_Y0D_hi_unq1),
    .out(Tile_X07_Y0D_hi_out)
);
mantle_wire__typeBit8 Tile_X07_Y0D_lo (
    .in(Tile_X07_Y0D_lo_unq1),
    .out(Tile_X07_Y0D_lo_out)
);
wire [15:0] Tile_X07_Y0D_tile_id_out;
assign Tile_X07_Y0D_tile_id_out = {Tile_X07_Y0D_lo_out[7],Tile_X07_Y0D_lo_out[7:6],Tile_X07_Y0D_lo_out[6:5],Tile_X07_Y0D_hi_out[5],Tile_X07_Y0D_hi_out[5:4],Tile_X07_Y0D_lo_out[3],Tile_X07_Y0D_lo_out[3:2],Tile_X07_Y0D_lo_out[2],Tile_X07_Y0D_hi_out[2:1],Tile_X07_Y0D_lo_out[0],Tile_X07_Y0D_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X07_Y0D_tile_id (
    .in(Tile_X07_Y0D_tile_id_in),
    .out(Tile_X07_Y0D_tile_id_out)
);
Tile_MemCore Tile_X07_Y0E (
    .SB_T0_EAST_SB_IN_B1(Tile_X08_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X08_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X07_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X07_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X07_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X07_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X07_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X07_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X07_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X07_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X07_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X07_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X06_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X06_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X07_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X07_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X08_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X08_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X07_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X07_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X07_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X07_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X07_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X07_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X07_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X07_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X07_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X07_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X06_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X06_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X07_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X07_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X08_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X08_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X07_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X07_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X07_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X07_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X07_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X07_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X07_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X07_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X07_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X07_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X06_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X06_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X07_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X07_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X08_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X08_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X07_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X07_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X07_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X07_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X07_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X07_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X07_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X07_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X07_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X07_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X06_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X06_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X07_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X07_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X08_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X08_Y0E_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X07_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X07_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X07_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X07_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X07_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X07_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X07_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X07_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X07_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X07_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X06_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X06_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X07_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X07_Y0E_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y0E_clk_pass_through_out_right),
    .clk_out(Tile_X07_Y0E_clk_out),
    .config_config_addr(Tile_X07_Y0D_config_out_config_addr),
    .config_config_data(Tile_X07_Y0D_config_out_config_data),
    .config_out_config_addr(Tile_X07_Y0E_config_out_config_addr),
    .config_out_config_data(Tile_X07_Y0E_config_out_config_data),
    .config_out_read(Tile_X07_Y0E_config_out_read),
    .config_out_write(Tile_X07_Y0E_config_out_write),
    .config_read(Tile_X07_Y0D_config_out_read),
    .config_write(Tile_X07_Y0D_config_out_write),
    .hi(Tile_X07_Y0E_hi_unq1),
    .lo(Tile_X07_Y0E_lo_unq1),
    .read_config_data(Tile_X07_Y0E_read_config_data),
    .read_config_data_in(Tile_X07_Y0D_read_config_data),
    .reset(Tile_X07_Y0D_reset_out),
    .reset_out(Tile_X07_Y0E_reset_out),
    .stall(Tile_X07_Y0D_stall_out),
    .stall_out(Tile_X07_Y0E_stall_out),
    .tile_id(Tile_X07_Y0E_tile_id_in)
);
mantle_wire__typeBit9 Tile_X07_Y0E_hi (
    .in(Tile_X07_Y0E_hi_unq1),
    .out(Tile_X07_Y0E_hi_out)
);
mantle_wire__typeBit8 Tile_X07_Y0E_lo (
    .in(Tile_X07_Y0E_lo_unq1),
    .out(Tile_X07_Y0E_lo_out)
);
wire [15:0] Tile_X07_Y0E_tile_id_out;
assign Tile_X07_Y0E_tile_id_out = {Tile_X07_Y0E_lo_out[7],Tile_X07_Y0E_lo_out[7:6],Tile_X07_Y0E_lo_out[6:5],Tile_X07_Y0E_hi_out[5],Tile_X07_Y0E_hi_out[5:4],Tile_X07_Y0E_lo_out[3],Tile_X07_Y0E_lo_out[3:2],Tile_X07_Y0E_lo_out[2],Tile_X07_Y0E_hi_out[2:1],Tile_X07_Y0E_hi_out[1],Tile_X07_Y0E_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X07_Y0E_tile_id (
    .in(Tile_X07_Y0E_tile_id_in),
    .out(Tile_X07_Y0E_tile_id_out)
);
Tile_MemCore Tile_X07_Y0F (
    .SB_T0_EAST_SB_IN_B1(Tile_X08_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X08_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X07_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X07_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X07_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X07_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X07_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X07_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X07_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X07_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X07_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X07_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X06_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X06_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X07_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X07_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X08_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X08_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X07_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X07_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X07_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X07_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X07_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X07_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X07_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X07_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X07_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X07_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X06_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X06_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X07_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X07_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X08_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X08_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X07_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X07_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X07_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X07_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X07_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X07_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X07_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X07_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X07_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X07_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X06_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X06_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X07_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X07_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X08_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X08_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X07_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X07_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X07_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X07_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X07_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X07_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X07_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X07_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X07_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X07_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X06_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X06_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X07_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X07_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X08_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X08_Y0F_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X07_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X07_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X07_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X07_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X07_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X07_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X07_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X07_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X07_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X07_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X06_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X06_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X07_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X07_Y0F_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y0F_clk_pass_through_out_right),
    .clk_out(Tile_X07_Y0F_clk_out),
    .config_config_addr(Tile_X07_Y0E_config_out_config_addr),
    .config_config_data(Tile_X07_Y0E_config_out_config_data),
    .config_out_config_addr(Tile_X07_Y0F_config_out_config_addr),
    .config_out_config_data(Tile_X07_Y0F_config_out_config_data),
    .config_out_read(Tile_X07_Y0F_config_out_read),
    .config_out_write(Tile_X07_Y0F_config_out_write),
    .config_read(Tile_X07_Y0E_config_out_read),
    .config_write(Tile_X07_Y0E_config_out_write),
    .hi(Tile_X07_Y0F_hi_unq1),
    .lo(Tile_X07_Y0F_lo_unq1),
    .read_config_data(Tile_X07_Y0F_read_config_data),
    .read_config_data_in(Tile_X07_Y0E_read_config_data),
    .reset(Tile_X07_Y0E_reset_out),
    .reset_out(Tile_X07_Y0F_reset_out),
    .stall(Tile_X07_Y0E_stall_out),
    .stall_out(Tile_X07_Y0F_stall_out),
    .tile_id(Tile_X07_Y0F_tile_id_in)
);
mantle_wire__typeBit9 Tile_X07_Y0F_hi (
    .in(Tile_X07_Y0F_hi_unq1),
    .out(Tile_X07_Y0F_hi_out)
);
mantle_wire__typeBit8 Tile_X07_Y0F_lo (
    .in(Tile_X07_Y0F_lo_unq1),
    .out(Tile_X07_Y0F_lo_out)
);
wire [15:0] Tile_X07_Y0F_tile_id_out;
assign Tile_X07_Y0F_tile_id_out = {Tile_X07_Y0F_lo_out[7],Tile_X07_Y0F_lo_out[7:6],Tile_X07_Y0F_lo_out[6:5],Tile_X07_Y0F_hi_out[5],Tile_X07_Y0F_hi_out[5:4],Tile_X07_Y0F_lo_out[3],Tile_X07_Y0F_lo_out[3:2],Tile_X07_Y0F_lo_out[2],Tile_X07_Y0F_hi_out[2:1],Tile_X07_Y0F_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X07_Y0F_tile_id (
    .in(Tile_X07_Y0F_tile_id_in),
    .out(Tile_X07_Y0F_tile_id_out)
);
Tile_MemCore Tile_X07_Y10 (
    .SB_T0_EAST_SB_IN_B1(Tile_X08_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X08_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X07_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X07_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X07_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X07_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X07_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X07_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T0_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X07_Y10_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X07_Y10_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X06_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X06_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X07_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X07_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X08_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X08_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X07_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X07_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X07_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X07_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X07_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X07_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T1_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X07_Y10_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X07_Y10_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X06_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X06_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X07_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X07_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X08_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X08_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X07_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X07_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X07_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X07_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X07_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X07_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T2_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X07_Y10_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X07_Y10_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X06_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X06_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X07_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X07_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X08_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X08_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X07_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X07_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X07_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X07_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X07_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X07_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T3_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X07_Y10_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X07_Y10_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X06_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X06_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X07_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X07_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X08_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X08_Y10_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X07_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X07_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X07_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X07_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X07_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X07_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T4_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X07_Y10_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X07_Y10_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X06_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X06_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X07_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X07_Y10_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X06_Y10_clk_pass_through_out_right),
    .clk_out(Tile_X07_Y10_clk_out),
    .config_config_addr(Tile_X07_Y0F_config_out_config_addr),
    .config_config_data(Tile_X07_Y0F_config_out_config_data),
    .config_out_config_addr(Tile_X07_Y10_config_out_config_addr),
    .config_out_config_data(Tile_X07_Y10_config_out_config_data),
    .config_out_read(Tile_X07_Y10_config_out_read),
    .config_out_write(Tile_X07_Y10_config_out_write),
    .config_read(Tile_X07_Y0F_config_out_read),
    .config_write(Tile_X07_Y0F_config_out_write),
    .hi(Tile_X07_Y10_hi_unq1),
    .lo(Tile_X07_Y10_lo_unq1),
    .read_config_data(Tile_X07_Y10_read_config_data),
    .read_config_data_in(Tile_X07_Y0F_read_config_data),
    .reset(Tile_X07_Y0F_reset_out),
    .reset_out(Tile_X07_Y10_reset_out),
    .stall(Tile_X07_Y0F_stall_out),
    .stall_out(Tile_X07_Y10_stall_out),
    .tile_id(Tile_X07_Y10_tile_id_in)
);
mantle_wire__typeBit9 Tile_X07_Y10_hi (
    .in(Tile_X07_Y10_hi_unq1),
    .out(Tile_X07_Y10_hi_out)
);
mantle_wire__typeBit8 Tile_X07_Y10_lo (
    .in(Tile_X07_Y10_lo_unq1),
    .out(Tile_X07_Y10_lo_out)
);
wire [15:0] Tile_X07_Y10_tile_id_out;
assign Tile_X07_Y10_tile_id_out = {Tile_X07_Y10_lo_out[7],Tile_X07_Y10_lo_out[7:6],Tile_X07_Y10_lo_out[6:5],Tile_X07_Y10_hi_out[5],Tile_X07_Y10_hi_out[5:4],Tile_X07_Y10_lo_out[3],Tile_X07_Y10_lo_out[3:2],Tile_X07_Y10_hi_out[2],Tile_X07_Y10_lo_out[1],Tile_X07_Y10_lo_out[1:0],Tile_X07_Y10_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X07_Y10_tile_id (
    .in(Tile_X07_Y10_tile_id_in),
    .out(Tile_X07_Y10_tile_id_out)
);
wire [15:0] Tile_X08_Y00_tile_id;
assign Tile_X08_Y00_tile_id = {Tile_X08_Y00_lo[7],Tile_X08_Y00_lo[7:6],Tile_X08_Y00_lo[6],Tile_X08_Y00_hi[6],Tile_X08_Y00_lo[5:4],Tile_X08_Y00_lo[4:3],Tile_X08_Y00_lo[3:2],Tile_X08_Y00_lo[2:1],Tile_X08_Y00_lo[1:0],Tile_X08_Y00_lo[0]};
Tile_io_core Tile_X08_Y00 (
    .tile_id(Tile_X08_Y00_tile_id),
    .glb2io_1(glb2io_1_X08_Y00),
    .f2io_1(Tile_X08_Y01_SB_T0_NORTH_SB_OUT_B1),
    .io2glb_1(Tile_X08_Y00_io2glb_1),
    .io2f_1(Tile_X08_Y00_io2f_1),
    .glb2io_16(glb2io_16_X08_Y00),
    .f2io_16(Tile_X08_Y01_SB_T0_NORTH_SB_OUT_B16),
    .io2glb_16(Tile_X08_Y00_io2glb_16),
    .io2f_16(Tile_X08_Y00_io2f_16),
    .hi(Tile_X08_Y00_hi),
    .lo(Tile_X08_Y00_lo)
);
Tile_PE Tile_X08_Y01 (
    .SB_T0_EAST_SB_IN_B1(Tile_X09_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X09_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X08_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X08_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X08_Y00_io2f_1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X08_Y00_io2f_16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X08_Y01_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X08_Y01_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X08_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X08_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X08_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X08_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X07_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X07_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X08_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X08_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X09_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X09_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X08_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X08_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X08_Y00_io2f_1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X08_Y00_io2f_16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X08_Y01_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X08_Y01_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X08_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X08_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X08_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X08_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X07_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X07_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X08_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X08_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X09_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X09_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X08_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X08_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X08_Y00_io2f_1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X08_Y00_io2f_16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X08_Y01_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X08_Y01_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X08_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X08_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X08_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X08_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X07_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X07_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X08_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X08_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X09_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X09_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X08_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X08_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X08_Y00_io2f_1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X08_Y00_io2f_16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X08_Y01_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X08_Y01_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X08_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X08_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X08_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X08_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X07_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X07_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X08_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X08_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X09_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X09_Y01_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X08_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X08_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X08_Y00_io2f_1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X08_Y00_io2f_16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X08_Y01_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X08_Y01_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X08_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X08_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X08_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X08_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X07_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X07_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X08_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X08_Y01_SB_T4_WEST_SB_OUT_B16),
    .clk(clk),
    .clk_out(Tile_X08_Y01_clk_out),
    .clk_pass_through(clk),
    .clk_pass_through_out_bot(Tile_X08_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X08_Y01_clk_pass_through_out_right),
    .config_config_addr(config_8_config_addr),
    .config_config_data(config_8_config_data),
    .config_out_config_addr(Tile_X08_Y01_config_out_config_addr),
    .config_out_config_data(Tile_X08_Y01_config_out_config_data),
    .config_out_read(Tile_X08_Y01_config_out_read),
    .config_out_write(Tile_X08_Y01_config_out_write),
    .config_read(config_8_read),
    .config_write(config_8_write),
    .hi(Tile_X08_Y01_hi),
    .lo(Tile_X08_Y01_lo_unq1),
    .read_config_data(Tile_X08_Y01_read_config_data),
    .read_config_data_in(const_0_32_out),
    .reset(reset),
    .reset_out(Tile_X08_Y01_reset_out),
    .stall(stall[8]),
    .stall_out(Tile_X08_Y01_stall_out),
    .tile_id(Tile_X08_Y01_tile_id_in)
);
mantle_wire__typeBit8 Tile_X08_Y01_lo (
    .in(Tile_X08_Y01_lo_unq1),
    .out(Tile_X08_Y01_lo_out)
);
wire [15:0] Tile_X08_Y01_tile_id_out;
assign Tile_X08_Y01_tile_id_out = {Tile_X08_Y01_lo_out[7],Tile_X08_Y01_lo_out[7:6],Tile_X08_Y01_lo_out[6],Tile_X08_Y01_hi[6],Tile_X08_Y01_lo_out[5:4],Tile_X08_Y01_lo_out[4:3],Tile_X08_Y01_lo_out[3:2],Tile_X08_Y01_lo_out[2:1],Tile_X08_Y01_lo_out[1:0],Tile_X08_Y01_hi[0]};
mantle_wire__typeBitIn16 Tile_X08_Y01_tile_id (
    .in(Tile_X08_Y01_tile_id_in),
    .out(Tile_X08_Y01_tile_id_out)
);
Tile_PE Tile_X08_Y02 (
    .SB_T0_EAST_SB_IN_B1(Tile_X09_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X09_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X08_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X08_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X08_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X08_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X08_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X08_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X08_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X08_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X08_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X08_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X07_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X07_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X08_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X08_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X09_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X09_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X08_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X08_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X08_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X08_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X08_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X08_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X08_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X08_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X08_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X08_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X07_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X07_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X08_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X08_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X09_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X09_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X08_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X08_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X08_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X08_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X08_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X08_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X08_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X08_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X08_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X08_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X07_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X07_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X08_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X08_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X09_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X09_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X08_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X08_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X08_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X08_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X08_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X08_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X08_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X08_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X08_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X08_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X07_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X07_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X08_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X08_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X09_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X09_Y02_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X08_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X08_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X08_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X08_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X08_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X08_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X08_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X08_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X08_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X08_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X07_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X07_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X08_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X08_Y02_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X08_Y01_clk_out),
    .clk_out(Tile_X08_Y02_clk_out),
    .clk_pass_through(Tile_X08_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X08_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X08_Y02_clk_pass_through_out_right),
    .config_config_addr(Tile_X08_Y01_config_out_config_addr),
    .config_config_data(Tile_X08_Y01_config_out_config_data),
    .config_out_config_addr(Tile_X08_Y02_config_out_config_addr),
    .config_out_config_data(Tile_X08_Y02_config_out_config_data),
    .config_out_read(Tile_X08_Y02_config_out_read),
    .config_out_write(Tile_X08_Y02_config_out_write),
    .config_read(Tile_X08_Y01_config_out_read),
    .config_write(Tile_X08_Y01_config_out_write),
    .hi(Tile_X08_Y02_hi),
    .lo(Tile_X08_Y02_lo_unq1),
    .read_config_data(Tile_X08_Y02_read_config_data),
    .read_config_data_in(Tile_X08_Y01_read_config_data),
    .reset(Tile_X08_Y01_reset_out),
    .reset_out(Tile_X08_Y02_reset_out),
    .stall(Tile_X08_Y01_stall_out),
    .stall_out(Tile_X08_Y02_stall_out),
    .tile_id(Tile_X08_Y02_tile_id_in)
);
mantle_wire__typeBit8 Tile_X08_Y02_lo (
    .in(Tile_X08_Y02_lo_unq1),
    .out(Tile_X08_Y02_lo_out)
);
wire [15:0] Tile_X08_Y02_tile_id_out;
assign Tile_X08_Y02_tile_id_out = {Tile_X08_Y02_lo_out[7],Tile_X08_Y02_lo_out[7:6],Tile_X08_Y02_lo_out[6],Tile_X08_Y02_hi[6],Tile_X08_Y02_lo_out[5:4],Tile_X08_Y02_lo_out[4:3],Tile_X08_Y02_lo_out[3:2],Tile_X08_Y02_lo_out[2:1],Tile_X08_Y02_lo_out[1],Tile_X08_Y02_hi[1],Tile_X08_Y02_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X08_Y02_tile_id (
    .in(Tile_X08_Y02_tile_id_in),
    .out(Tile_X08_Y02_tile_id_out)
);
Tile_PE Tile_X08_Y03 (
    .SB_T0_EAST_SB_IN_B1(Tile_X09_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X09_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X08_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X08_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X08_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X08_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X08_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X08_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X08_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X08_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X08_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X08_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X07_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X07_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X08_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X08_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X09_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X09_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X08_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X08_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X08_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X08_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X08_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X08_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X08_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X08_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X08_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X08_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X07_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X07_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X08_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X08_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X09_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X09_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X08_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X08_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X08_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X08_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X08_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X08_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X08_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X08_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X08_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X08_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X07_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X07_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X08_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X08_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X09_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X09_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X08_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X08_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X08_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X08_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X08_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X08_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X08_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X08_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X08_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X08_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X07_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X07_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X08_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X08_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X09_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X09_Y03_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X08_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X08_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X08_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X08_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X08_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X08_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X08_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X08_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X08_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X08_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X07_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X07_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X08_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X08_Y03_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X08_Y02_clk_out),
    .clk_out(Tile_X08_Y03_clk_out),
    .clk_pass_through(Tile_X08_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X08_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X08_Y03_clk_pass_through_out_right),
    .config_config_addr(Tile_X08_Y02_config_out_config_addr),
    .config_config_data(Tile_X08_Y02_config_out_config_data),
    .config_out_config_addr(Tile_X08_Y03_config_out_config_addr),
    .config_out_config_data(Tile_X08_Y03_config_out_config_data),
    .config_out_read(Tile_X08_Y03_config_out_read),
    .config_out_write(Tile_X08_Y03_config_out_write),
    .config_read(Tile_X08_Y02_config_out_read),
    .config_write(Tile_X08_Y02_config_out_write),
    .hi(Tile_X08_Y03_hi_unq1),
    .lo(Tile_X08_Y03_lo_unq1),
    .read_config_data(Tile_X08_Y03_read_config_data),
    .read_config_data_in(Tile_X08_Y02_read_config_data),
    .reset(Tile_X08_Y02_reset_out),
    .reset_out(Tile_X08_Y03_reset_out),
    .stall(Tile_X08_Y02_stall_out),
    .stall_out(Tile_X08_Y03_stall_out),
    .tile_id(Tile_X08_Y03_tile_id_in)
);
mantle_wire__typeBit9 Tile_X08_Y03_hi (
    .in(Tile_X08_Y03_hi_unq1),
    .out(Tile_X08_Y03_hi_out)
);
mantle_wire__typeBit8 Tile_X08_Y03_lo (
    .in(Tile_X08_Y03_lo_unq1),
    .out(Tile_X08_Y03_lo_out)
);
wire [15:0] Tile_X08_Y03_tile_id_out;
assign Tile_X08_Y03_tile_id_out = {Tile_X08_Y03_lo_out[7],Tile_X08_Y03_lo_out[7:6],Tile_X08_Y03_lo_out[6],Tile_X08_Y03_hi_out[6],Tile_X08_Y03_lo_out[5:4],Tile_X08_Y03_lo_out[4:3],Tile_X08_Y03_lo_out[3:2],Tile_X08_Y03_lo_out[2:1],Tile_X08_Y03_lo_out[1],Tile_X08_Y03_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X08_Y03_tile_id (
    .in(Tile_X08_Y03_tile_id_in),
    .out(Tile_X08_Y03_tile_id_out)
);
Tile_PE Tile_X08_Y04 (
    .SB_T0_EAST_SB_IN_B1(Tile_X09_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X09_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X08_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X08_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X08_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X08_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X08_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X08_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X08_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X08_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X08_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X08_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X07_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X07_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X08_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X08_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X09_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X09_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X08_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X08_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X08_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X08_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X08_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X08_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X08_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X08_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X08_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X08_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X07_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X07_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X08_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X08_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X09_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X09_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X08_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X08_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X08_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X08_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X08_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X08_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X08_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X08_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X08_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X08_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X07_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X07_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X08_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X08_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X09_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X09_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X08_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X08_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X08_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X08_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X08_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X08_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X08_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X08_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X08_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X08_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X07_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X07_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X08_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X08_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X09_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X09_Y04_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X08_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X08_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X08_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X08_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X08_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X08_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X08_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X08_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X08_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X08_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X07_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X07_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X08_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X08_Y04_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X08_Y03_clk_out),
    .clk_out(Tile_X08_Y04_clk_out),
    .clk_pass_through(Tile_X08_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X08_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X08_Y04_clk_pass_through_out_right),
    .config_config_addr(Tile_X08_Y03_config_out_config_addr),
    .config_config_data(Tile_X08_Y03_config_out_config_data),
    .config_out_config_addr(Tile_X08_Y04_config_out_config_addr),
    .config_out_config_data(Tile_X08_Y04_config_out_config_data),
    .config_out_read(Tile_X08_Y04_config_out_read),
    .config_out_write(Tile_X08_Y04_config_out_write),
    .config_read(Tile_X08_Y03_config_out_read),
    .config_write(Tile_X08_Y03_config_out_write),
    .hi(Tile_X08_Y04_hi),
    .lo(Tile_X08_Y04_lo_unq1),
    .read_config_data(Tile_X08_Y04_read_config_data),
    .read_config_data_in(Tile_X08_Y03_read_config_data),
    .reset(Tile_X08_Y03_reset_out),
    .reset_out(Tile_X08_Y04_reset_out),
    .stall(Tile_X08_Y03_stall_out),
    .stall_out(Tile_X08_Y04_stall_out),
    .tile_id(Tile_X08_Y04_tile_id_in)
);
mantle_wire__typeBit8 Tile_X08_Y04_lo (
    .in(Tile_X08_Y04_lo_unq1),
    .out(Tile_X08_Y04_lo_out)
);
wire [15:0] Tile_X08_Y04_tile_id_out;
assign Tile_X08_Y04_tile_id_out = {Tile_X08_Y04_lo_out[7],Tile_X08_Y04_lo_out[7:6],Tile_X08_Y04_lo_out[6],Tile_X08_Y04_hi[6],Tile_X08_Y04_lo_out[5:4],Tile_X08_Y04_lo_out[4:3],Tile_X08_Y04_lo_out[3:2],Tile_X08_Y04_lo_out[2:1],Tile_X08_Y04_hi[1],Tile_X08_Y04_lo_out[0],Tile_X08_Y04_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X08_Y04_tile_id (
    .in(Tile_X08_Y04_tile_id_in),
    .out(Tile_X08_Y04_tile_id_out)
);
Tile_PE Tile_X08_Y05 (
    .SB_T0_EAST_SB_IN_B1(Tile_X09_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X09_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X08_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X08_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X08_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X08_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X08_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X08_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X08_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X08_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X08_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X08_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X07_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X07_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X08_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X08_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X09_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X09_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X08_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X08_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X08_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X08_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X08_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X08_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X08_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X08_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X08_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X08_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X07_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X07_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X08_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X08_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X09_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X09_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X08_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X08_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X08_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X08_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X08_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X08_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X08_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X08_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X08_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X08_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X07_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X07_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X08_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X08_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X09_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X09_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X08_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X08_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X08_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X08_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X08_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X08_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X08_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X08_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X08_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X08_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X07_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X07_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X08_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X08_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X09_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X09_Y05_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X08_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X08_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X08_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X08_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X08_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X08_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X08_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X08_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X08_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X08_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X07_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X07_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X08_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X08_Y05_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X08_Y04_clk_out),
    .clk_out(Tile_X08_Y05_clk_out),
    .clk_pass_through(Tile_X08_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X08_Y05_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X08_Y05_clk_pass_through_out_right),
    .config_config_addr(Tile_X08_Y04_config_out_config_addr),
    .config_config_data(Tile_X08_Y04_config_out_config_data),
    .config_out_config_addr(Tile_X08_Y05_config_out_config_addr),
    .config_out_config_data(Tile_X08_Y05_config_out_config_data),
    .config_out_read(Tile_X08_Y05_config_out_read),
    .config_out_write(Tile_X08_Y05_config_out_write),
    .config_read(Tile_X08_Y04_config_out_read),
    .config_write(Tile_X08_Y04_config_out_write),
    .hi(Tile_X08_Y05_hi),
    .lo(Tile_X08_Y05_lo_unq1),
    .read_config_data(Tile_X08_Y05_read_config_data),
    .read_config_data_in(Tile_X08_Y04_read_config_data),
    .reset(Tile_X08_Y04_reset_out),
    .reset_out(Tile_X08_Y05_reset_out),
    .stall(Tile_X08_Y04_stall_out),
    .stall_out(Tile_X08_Y05_stall_out),
    .tile_id(Tile_X08_Y05_tile_id_in)
);
mantle_wire__typeBit8 Tile_X08_Y05_lo (
    .in(Tile_X08_Y05_lo_unq1),
    .out(Tile_X08_Y05_lo_out)
);
wire [15:0] Tile_X08_Y05_tile_id_out;
assign Tile_X08_Y05_tile_id_out = {Tile_X08_Y05_lo_out[7],Tile_X08_Y05_lo_out[7:6],Tile_X08_Y05_lo_out[6],Tile_X08_Y05_hi[6],Tile_X08_Y05_lo_out[5:4],Tile_X08_Y05_lo_out[4:3],Tile_X08_Y05_lo_out[3:2],Tile_X08_Y05_lo_out[2:1],Tile_X08_Y05_hi[1],Tile_X08_Y05_lo_out[0],Tile_X08_Y05_hi[0]};
mantle_wire__typeBitIn16 Tile_X08_Y05_tile_id (
    .in(Tile_X08_Y05_tile_id_in),
    .out(Tile_X08_Y05_tile_id_out)
);
Tile_PE Tile_X08_Y06 (
    .SB_T0_EAST_SB_IN_B1(Tile_X09_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X09_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X08_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X08_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X08_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X08_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X08_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X08_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X08_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X08_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X08_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X08_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X07_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X07_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X08_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X08_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X09_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X09_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X08_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X08_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X08_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X08_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X08_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X08_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X08_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X08_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X08_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X08_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X07_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X07_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X08_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X08_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X09_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X09_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X08_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X08_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X08_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X08_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X08_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X08_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X08_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X08_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X08_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X08_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X07_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X07_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X08_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X08_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X09_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X09_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X08_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X08_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X08_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X08_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X08_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X08_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X08_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X08_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X08_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X08_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X07_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X07_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X08_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X08_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X09_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X09_Y06_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X08_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X08_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X08_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X08_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X08_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X08_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X08_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X08_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X08_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X08_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X07_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X07_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X08_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X08_Y06_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X08_Y05_clk_out),
    .clk_out(Tile_X08_Y06_clk_out),
    .clk_pass_through(Tile_X08_Y05_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X08_Y06_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X08_Y06_clk_pass_through_out_right),
    .config_config_addr(Tile_X08_Y05_config_out_config_addr),
    .config_config_data(Tile_X08_Y05_config_out_config_data),
    .config_out_config_addr(Tile_X08_Y06_config_out_config_addr),
    .config_out_config_data(Tile_X08_Y06_config_out_config_data),
    .config_out_read(Tile_X08_Y06_config_out_read),
    .config_out_write(Tile_X08_Y06_config_out_write),
    .config_read(Tile_X08_Y05_config_out_read),
    .config_write(Tile_X08_Y05_config_out_write),
    .hi(Tile_X08_Y06_hi),
    .lo(Tile_X08_Y06_lo_unq1),
    .read_config_data(Tile_X08_Y06_read_config_data),
    .read_config_data_in(Tile_X08_Y05_read_config_data),
    .reset(Tile_X08_Y05_reset_out),
    .reset_out(Tile_X08_Y06_reset_out),
    .stall(Tile_X08_Y05_stall_out),
    .stall_out(Tile_X08_Y06_stall_out),
    .tile_id(Tile_X08_Y06_tile_id_in)
);
mantle_wire__typeBit8 Tile_X08_Y06_lo (
    .in(Tile_X08_Y06_lo_unq1),
    .out(Tile_X08_Y06_lo_out)
);
wire [15:0] Tile_X08_Y06_tile_id_out;
assign Tile_X08_Y06_tile_id_out = {Tile_X08_Y06_lo_out[7],Tile_X08_Y06_lo_out[7:6],Tile_X08_Y06_lo_out[6],Tile_X08_Y06_hi[6],Tile_X08_Y06_lo_out[5:4],Tile_X08_Y06_lo_out[4:3],Tile_X08_Y06_lo_out[3:2],Tile_X08_Y06_lo_out[2:1],Tile_X08_Y06_hi[1],Tile_X08_Y06_hi[1],Tile_X08_Y06_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X08_Y06_tile_id (
    .in(Tile_X08_Y06_tile_id_in),
    .out(Tile_X08_Y06_tile_id_out)
);
Tile_PE Tile_X08_Y07 (
    .SB_T0_EAST_SB_IN_B1(Tile_X09_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X09_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X08_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X08_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X08_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X08_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X08_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X08_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X08_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X08_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X08_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X08_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X07_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X07_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X08_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X08_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X09_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X09_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X08_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X08_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X08_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X08_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X08_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X08_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X08_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X08_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X08_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X08_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X07_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X07_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X08_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X08_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X09_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X09_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X08_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X08_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X08_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X08_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X08_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X08_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X08_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X08_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X08_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X08_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X07_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X07_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X08_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X08_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X09_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X09_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X08_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X08_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X08_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X08_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X08_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X08_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X08_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X08_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X08_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X08_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X07_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X07_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X08_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X08_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X09_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X09_Y07_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X08_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X08_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X08_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X08_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X08_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X08_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X08_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X08_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X08_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X08_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X07_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X07_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X08_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X08_Y07_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X08_Y06_clk_out),
    .clk_out(Tile_X08_Y07_clk_out),
    .clk_pass_through(Tile_X08_Y06_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X08_Y07_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X08_Y07_clk_pass_through_out_right),
    .config_config_addr(Tile_X08_Y06_config_out_config_addr),
    .config_config_data(Tile_X08_Y06_config_out_config_data),
    .config_out_config_addr(Tile_X08_Y07_config_out_config_addr),
    .config_out_config_data(Tile_X08_Y07_config_out_config_data),
    .config_out_read(Tile_X08_Y07_config_out_read),
    .config_out_write(Tile_X08_Y07_config_out_write),
    .config_read(Tile_X08_Y06_config_out_read),
    .config_write(Tile_X08_Y06_config_out_write),
    .hi(Tile_X08_Y07_hi_unq1),
    .lo(Tile_X08_Y07_lo_unq1),
    .read_config_data(Tile_X08_Y07_read_config_data),
    .read_config_data_in(Tile_X08_Y06_read_config_data),
    .reset(Tile_X08_Y06_reset_out),
    .reset_out(Tile_X08_Y07_reset_out),
    .stall(Tile_X08_Y06_stall_out),
    .stall_out(Tile_X08_Y07_stall_out),
    .tile_id(Tile_X08_Y07_tile_id_in)
);
mantle_wire__typeBit9 Tile_X08_Y07_hi (
    .in(Tile_X08_Y07_hi_unq1),
    .out(Tile_X08_Y07_hi_out)
);
mantle_wire__typeBit8 Tile_X08_Y07_lo (
    .in(Tile_X08_Y07_lo_unq1),
    .out(Tile_X08_Y07_lo_out)
);
wire [15:0] Tile_X08_Y07_tile_id_out;
assign Tile_X08_Y07_tile_id_out = {Tile_X08_Y07_lo_out[7],Tile_X08_Y07_lo_out[7:6],Tile_X08_Y07_lo_out[6],Tile_X08_Y07_hi_out[6],Tile_X08_Y07_lo_out[5:4],Tile_X08_Y07_lo_out[4:3],Tile_X08_Y07_lo_out[3:2],Tile_X08_Y07_lo_out[2:1],Tile_X08_Y07_hi_out[1],Tile_X08_Y07_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X08_Y07_tile_id (
    .in(Tile_X08_Y07_tile_id_in),
    .out(Tile_X08_Y07_tile_id_out)
);
Tile_PE Tile_X08_Y08 (
    .SB_T0_EAST_SB_IN_B1(Tile_X09_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X09_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X08_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X08_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X08_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X08_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X08_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X08_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X08_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X08_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X08_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X08_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X07_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X07_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X08_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X08_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X09_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X09_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X08_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X08_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X08_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X08_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X08_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X08_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X08_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X08_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X08_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X08_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X07_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X07_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X08_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X08_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X09_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X09_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X08_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X08_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X08_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X08_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X08_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X08_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X08_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X08_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X08_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X08_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X07_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X07_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X08_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X08_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X09_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X09_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X08_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X08_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X08_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X08_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X08_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X08_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X08_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X08_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X08_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X08_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X07_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X07_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X08_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X08_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X09_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X09_Y08_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X08_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X08_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X08_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X08_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X08_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X08_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X08_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X08_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X08_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X08_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X07_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X07_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X08_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X08_Y08_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X08_Y07_clk_out),
    .clk_out(Tile_X08_Y08_clk_out),
    .clk_pass_through(Tile_X08_Y07_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X08_Y08_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X08_Y08_clk_pass_through_out_right),
    .config_config_addr(Tile_X08_Y07_config_out_config_addr),
    .config_config_data(Tile_X08_Y07_config_out_config_data),
    .config_out_config_addr(Tile_X08_Y08_config_out_config_addr),
    .config_out_config_data(Tile_X08_Y08_config_out_config_data),
    .config_out_read(Tile_X08_Y08_config_out_read),
    .config_out_write(Tile_X08_Y08_config_out_write),
    .config_read(Tile_X08_Y07_config_out_read),
    .config_write(Tile_X08_Y07_config_out_write),
    .hi(Tile_X08_Y08_hi),
    .lo(Tile_X08_Y08_lo_unq1),
    .read_config_data(Tile_X08_Y08_read_config_data),
    .read_config_data_in(Tile_X08_Y07_read_config_data),
    .reset(Tile_X08_Y07_reset_out),
    .reset_out(Tile_X08_Y08_reset_out),
    .stall(Tile_X08_Y07_stall_out),
    .stall_out(Tile_X08_Y08_stall_out),
    .tile_id(Tile_X08_Y08_tile_id_in)
);
mantle_wire__typeBit8 Tile_X08_Y08_lo (
    .in(Tile_X08_Y08_lo_unq1),
    .out(Tile_X08_Y08_lo_out)
);
wire [15:0] Tile_X08_Y08_tile_id_out;
assign Tile_X08_Y08_tile_id_out = {Tile_X08_Y08_lo_out[7],Tile_X08_Y08_lo_out[7:6],Tile_X08_Y08_lo_out[6],Tile_X08_Y08_hi[6],Tile_X08_Y08_lo_out[5:4],Tile_X08_Y08_lo_out[4:3],Tile_X08_Y08_lo_out[3:2],Tile_X08_Y08_lo_out[2],Tile_X08_Y08_hi[2],Tile_X08_Y08_lo_out[1:0],Tile_X08_Y08_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X08_Y08_tile_id (
    .in(Tile_X08_Y08_tile_id_in),
    .out(Tile_X08_Y08_tile_id_out)
);
Tile_PE Tile_X08_Y09 (
    .SB_T0_EAST_SB_IN_B1(Tile_X09_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X09_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X08_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X08_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X08_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X08_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X08_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X08_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X08_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X08_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X08_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X08_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X07_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X07_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X08_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X08_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X09_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X09_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X08_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X08_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X08_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X08_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X08_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X08_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X08_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X08_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X08_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X08_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X07_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X07_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X08_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X08_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X09_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X09_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X08_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X08_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X08_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X08_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X08_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X08_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X08_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X08_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X08_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X08_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X07_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X07_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X08_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X08_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X09_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X09_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X08_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X08_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X08_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X08_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X08_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X08_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X08_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X08_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X08_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X08_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X07_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X07_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X08_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X08_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X09_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X09_Y09_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X08_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X08_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X08_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X08_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X08_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X08_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X08_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X08_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X08_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X08_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X07_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X07_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X08_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X08_Y09_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X08_Y08_clk_out),
    .clk_out(Tile_X08_Y09_clk_out),
    .clk_pass_through(Tile_X08_Y08_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X08_Y09_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X08_Y09_clk_pass_through_out_right),
    .config_config_addr(ConfigPipeStage_inst8_config_out_config_addr),
    .config_config_data(ConfigPipeStage_inst8_config_out_config_data),
    .config_out_config_addr(Tile_X08_Y09_config_out_config_addr),
    .config_out_config_data(Tile_X08_Y09_config_out_config_data),
    .config_out_read(Tile_X08_Y09_config_out_read),
    .config_out_write(Tile_X08_Y09_config_out_write),
    .config_read(ConfigPipeStage_inst8_config_out_read),
    .config_write(ConfigPipeStage_inst8_config_out_write),
    .hi(Tile_X08_Y09_hi),
    .lo(Tile_X08_Y09_lo_unq1),
    .read_config_data(Tile_X08_Y09_read_config_data),
    .read_config_data_in(Tile_X08_Y08_read_config_data),
    .reset(Tile_X08_Y08_reset_out),
    .reset_out(Tile_X08_Y09_reset_out),
    .stall(Tile_X08_Y08_stall_out),
    .stall_out(Tile_X08_Y09_stall_out),
    .tile_id(Tile_X08_Y09_tile_id_in)
);
mantle_wire__typeBit8 Tile_X08_Y09_lo (
    .in(Tile_X08_Y09_lo_unq1),
    .out(Tile_X08_Y09_lo_out)
);
wire [15:0] Tile_X08_Y09_tile_id_out;
assign Tile_X08_Y09_tile_id_out = {Tile_X08_Y09_lo_out[7],Tile_X08_Y09_lo_out[7:6],Tile_X08_Y09_lo_out[6],Tile_X08_Y09_hi[6],Tile_X08_Y09_lo_out[5:4],Tile_X08_Y09_lo_out[4:3],Tile_X08_Y09_lo_out[3:2],Tile_X08_Y09_lo_out[2],Tile_X08_Y09_hi[2],Tile_X08_Y09_lo_out[1:0],Tile_X08_Y09_hi[0]};
mantle_wire__typeBitIn16 Tile_X08_Y09_tile_id (
    .in(Tile_X08_Y09_tile_id_in),
    .out(Tile_X08_Y09_tile_id_out)
);
Tile_PE Tile_X08_Y0A (
    .SB_T0_EAST_SB_IN_B1(Tile_X09_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X09_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X08_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X08_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X08_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X08_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X08_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X08_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X08_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X08_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X08_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X08_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X07_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X07_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X08_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X08_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X09_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X09_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X08_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X08_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X08_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X08_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X08_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X08_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X08_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X08_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X08_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X08_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X07_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X07_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X08_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X08_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X09_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X09_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X08_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X08_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X08_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X08_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X08_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X08_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X08_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X08_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X08_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X08_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X07_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X07_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X08_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X08_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X09_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X09_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X08_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X08_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X08_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X08_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X08_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X08_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X08_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X08_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X08_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X08_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X07_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X07_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X08_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X08_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X09_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X09_Y0A_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X08_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X08_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X08_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X08_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X08_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X08_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X08_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X08_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X08_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X08_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X07_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X07_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X08_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X08_Y0A_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X08_Y09_clk_out),
    .clk_out(Tile_X08_Y0A_clk_out),
    .clk_pass_through(Tile_X08_Y09_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X08_Y0A_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X08_Y0A_clk_pass_through_out_right),
    .config_config_addr(Tile_X08_Y09_config_out_config_addr),
    .config_config_data(Tile_X08_Y09_config_out_config_data),
    .config_out_config_addr(Tile_X08_Y0A_config_out_config_addr),
    .config_out_config_data(Tile_X08_Y0A_config_out_config_data),
    .config_out_read(Tile_X08_Y0A_config_out_read),
    .config_out_write(Tile_X08_Y0A_config_out_write),
    .config_read(Tile_X08_Y09_config_out_read),
    .config_write(Tile_X08_Y09_config_out_write),
    .hi(Tile_X08_Y0A_hi),
    .lo(Tile_X08_Y0A_lo_unq1),
    .read_config_data(Tile_X08_Y0A_read_config_data),
    .read_config_data_in(Tile_X08_Y09_read_config_data),
    .reset(Tile_X08_Y09_reset_out),
    .reset_out(Tile_X08_Y0A_reset_out),
    .stall(Tile_X08_Y09_stall_out),
    .stall_out(Tile_X08_Y0A_stall_out),
    .tile_id(Tile_X08_Y0A_tile_id_in)
);
mantle_wire__typeBit8 Tile_X08_Y0A_lo (
    .in(Tile_X08_Y0A_lo_unq1),
    .out(Tile_X08_Y0A_lo_out)
);
wire [15:0] Tile_X08_Y0A_tile_id_out;
assign Tile_X08_Y0A_tile_id_out = {Tile_X08_Y0A_lo_out[7],Tile_X08_Y0A_lo_out[7:6],Tile_X08_Y0A_lo_out[6],Tile_X08_Y0A_hi[6],Tile_X08_Y0A_lo_out[5:4],Tile_X08_Y0A_lo_out[4:3],Tile_X08_Y0A_lo_out[3:2],Tile_X08_Y0A_lo_out[2],Tile_X08_Y0A_hi[2],Tile_X08_Y0A_lo_out[1],Tile_X08_Y0A_hi[1],Tile_X08_Y0A_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X08_Y0A_tile_id (
    .in(Tile_X08_Y0A_tile_id_in),
    .out(Tile_X08_Y0A_tile_id_out)
);
Tile_PE Tile_X08_Y0B (
    .SB_T0_EAST_SB_IN_B1(Tile_X09_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X09_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X08_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X08_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X08_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X08_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X08_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X08_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X08_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X08_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X08_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X08_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X07_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X07_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X08_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X08_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X09_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X09_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X08_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X08_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X08_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X08_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X08_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X08_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X08_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X08_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X08_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X08_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X07_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X07_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X08_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X08_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X09_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X09_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X08_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X08_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X08_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X08_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X08_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X08_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X08_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X08_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X08_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X08_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X07_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X07_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X08_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X08_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X09_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X09_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X08_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X08_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X08_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X08_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X08_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X08_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X08_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X08_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X08_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X08_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X07_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X07_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X08_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X08_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X09_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X09_Y0B_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X08_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X08_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X08_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X08_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X08_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X08_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X08_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X08_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X08_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X08_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X07_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X07_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X08_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X08_Y0B_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X08_Y0A_clk_out),
    .clk_out(Tile_X08_Y0B_clk_out),
    .clk_pass_through(Tile_X08_Y0A_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X08_Y0B_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X08_Y0B_clk_pass_through_out_right),
    .config_config_addr(Tile_X08_Y0A_config_out_config_addr),
    .config_config_data(Tile_X08_Y0A_config_out_config_data),
    .config_out_config_addr(Tile_X08_Y0B_config_out_config_addr),
    .config_out_config_data(Tile_X08_Y0B_config_out_config_data),
    .config_out_read(Tile_X08_Y0B_config_out_read),
    .config_out_write(Tile_X08_Y0B_config_out_write),
    .config_read(Tile_X08_Y0A_config_out_read),
    .config_write(Tile_X08_Y0A_config_out_write),
    .hi(Tile_X08_Y0B_hi_unq1),
    .lo(Tile_X08_Y0B_lo_unq1),
    .read_config_data(Tile_X08_Y0B_read_config_data),
    .read_config_data_in(Tile_X08_Y0A_read_config_data),
    .reset(Tile_X08_Y0A_reset_out),
    .reset_out(Tile_X08_Y0B_reset_out),
    .stall(Tile_X08_Y0A_stall_out),
    .stall_out(Tile_X08_Y0B_stall_out),
    .tile_id(Tile_X08_Y0B_tile_id_in)
);
mantle_wire__typeBit9 Tile_X08_Y0B_hi (
    .in(Tile_X08_Y0B_hi_unq1),
    .out(Tile_X08_Y0B_hi_out)
);
mantle_wire__typeBit8 Tile_X08_Y0B_lo (
    .in(Tile_X08_Y0B_lo_unq1),
    .out(Tile_X08_Y0B_lo_out)
);
wire [15:0] Tile_X08_Y0B_tile_id_out;
assign Tile_X08_Y0B_tile_id_out = {Tile_X08_Y0B_lo_out[7],Tile_X08_Y0B_lo_out[7:6],Tile_X08_Y0B_lo_out[6],Tile_X08_Y0B_hi_out[6],Tile_X08_Y0B_lo_out[5:4],Tile_X08_Y0B_lo_out[4:3],Tile_X08_Y0B_lo_out[3:2],Tile_X08_Y0B_lo_out[2],Tile_X08_Y0B_hi_out[2],Tile_X08_Y0B_lo_out[1],Tile_X08_Y0B_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X08_Y0B_tile_id (
    .in(Tile_X08_Y0B_tile_id_in),
    .out(Tile_X08_Y0B_tile_id_out)
);
Tile_PE Tile_X08_Y0C (
    .SB_T0_EAST_SB_IN_B1(Tile_X09_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X09_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X08_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X08_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X08_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X08_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X08_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X08_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X08_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X08_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X08_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X08_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X07_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X07_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X08_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X08_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X09_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X09_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X08_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X08_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X08_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X08_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X08_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X08_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X08_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X08_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X08_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X08_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X07_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X07_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X08_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X08_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X09_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X09_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X08_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X08_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X08_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X08_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X08_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X08_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X08_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X08_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X08_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X08_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X07_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X07_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X08_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X08_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X09_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X09_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X08_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X08_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X08_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X08_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X08_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X08_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X08_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X08_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X08_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X08_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X07_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X07_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X08_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X08_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X09_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X09_Y0C_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X08_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X08_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X08_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X08_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X08_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X08_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X08_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X08_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X08_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X08_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X07_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X07_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X08_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X08_Y0C_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X08_Y0B_clk_out),
    .clk_out(Tile_X08_Y0C_clk_out),
    .clk_pass_through(Tile_X08_Y0B_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X08_Y0C_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X08_Y0C_clk_pass_through_out_right),
    .config_config_addr(Tile_X08_Y0B_config_out_config_addr),
    .config_config_data(Tile_X08_Y0B_config_out_config_data),
    .config_out_config_addr(Tile_X08_Y0C_config_out_config_addr),
    .config_out_config_data(Tile_X08_Y0C_config_out_config_data),
    .config_out_read(Tile_X08_Y0C_config_out_read),
    .config_out_write(Tile_X08_Y0C_config_out_write),
    .config_read(Tile_X08_Y0B_config_out_read),
    .config_write(Tile_X08_Y0B_config_out_write),
    .hi(Tile_X08_Y0C_hi_unq1),
    .lo(Tile_X08_Y0C_lo_unq1),
    .read_config_data(Tile_X08_Y0C_read_config_data),
    .read_config_data_in(Tile_X08_Y0B_read_config_data),
    .reset(Tile_X08_Y0B_reset_out),
    .reset_out(Tile_X08_Y0C_reset_out),
    .stall(Tile_X08_Y0B_stall_out),
    .stall_out(Tile_X08_Y0C_stall_out),
    .tile_id(Tile_X08_Y0C_tile_id_in)
);
mantle_wire__typeBit9 Tile_X08_Y0C_hi (
    .in(Tile_X08_Y0C_hi_unq1),
    .out(Tile_X08_Y0C_hi_out)
);
mantle_wire__typeBit8 Tile_X08_Y0C_lo (
    .in(Tile_X08_Y0C_lo_unq1),
    .out(Tile_X08_Y0C_lo_out)
);
wire [15:0] Tile_X08_Y0C_tile_id_out;
assign Tile_X08_Y0C_tile_id_out = {Tile_X08_Y0C_lo_out[7],Tile_X08_Y0C_lo_out[7:6],Tile_X08_Y0C_lo_out[6],Tile_X08_Y0C_hi_out[6],Tile_X08_Y0C_lo_out[5:4],Tile_X08_Y0C_lo_out[4:3],Tile_X08_Y0C_lo_out[3:2],Tile_X08_Y0C_lo_out[2],Tile_X08_Y0C_hi_out[2:1],Tile_X08_Y0C_lo_out[0],Tile_X08_Y0C_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X08_Y0C_tile_id (
    .in(Tile_X08_Y0C_tile_id_in),
    .out(Tile_X08_Y0C_tile_id_out)
);
Tile_PE Tile_X08_Y0D (
    .SB_T0_EAST_SB_IN_B1(Tile_X09_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X09_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X08_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X08_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X08_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X08_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X08_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X08_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X08_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X08_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X08_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X08_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X07_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X07_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X08_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X08_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X09_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X09_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X08_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X08_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X08_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X08_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X08_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X08_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X08_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X08_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X08_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X08_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X07_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X07_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X08_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X08_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X09_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X09_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X08_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X08_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X08_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X08_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X08_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X08_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X08_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X08_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X08_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X08_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X07_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X07_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X08_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X08_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X09_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X09_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X08_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X08_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X08_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X08_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X08_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X08_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X08_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X08_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X08_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X08_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X07_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X07_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X08_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X08_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X09_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X09_Y0D_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X08_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X08_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X08_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X08_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X08_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X08_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X08_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X08_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X08_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X08_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X07_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X07_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X08_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X08_Y0D_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X08_Y0C_clk_out),
    .clk_out(Tile_X08_Y0D_clk_out),
    .clk_pass_through(Tile_X08_Y0C_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X08_Y0D_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X08_Y0D_clk_pass_through_out_right),
    .config_config_addr(Tile_X08_Y0C_config_out_config_addr),
    .config_config_data(Tile_X08_Y0C_config_out_config_data),
    .config_out_config_addr(Tile_X08_Y0D_config_out_config_addr),
    .config_out_config_data(Tile_X08_Y0D_config_out_config_data),
    .config_out_read(Tile_X08_Y0D_config_out_read),
    .config_out_write(Tile_X08_Y0D_config_out_write),
    .config_read(Tile_X08_Y0C_config_out_read),
    .config_write(Tile_X08_Y0C_config_out_write),
    .hi(Tile_X08_Y0D_hi_unq1),
    .lo(Tile_X08_Y0D_lo_unq1),
    .read_config_data(Tile_X08_Y0D_read_config_data),
    .read_config_data_in(Tile_X08_Y0C_read_config_data),
    .reset(Tile_X08_Y0C_reset_out),
    .reset_out(Tile_X08_Y0D_reset_out),
    .stall(Tile_X08_Y0C_stall_out),
    .stall_out(Tile_X08_Y0D_stall_out),
    .tile_id(Tile_X08_Y0D_tile_id_in)
);
mantle_wire__typeBit9 Tile_X08_Y0D_hi (
    .in(Tile_X08_Y0D_hi_unq1),
    .out(Tile_X08_Y0D_hi_out)
);
mantle_wire__typeBit8 Tile_X08_Y0D_lo (
    .in(Tile_X08_Y0D_lo_unq1),
    .out(Tile_X08_Y0D_lo_out)
);
wire [15:0] Tile_X08_Y0D_tile_id_out;
assign Tile_X08_Y0D_tile_id_out = {Tile_X08_Y0D_lo_out[7],Tile_X08_Y0D_lo_out[7:6],Tile_X08_Y0D_lo_out[6],Tile_X08_Y0D_hi_out[6],Tile_X08_Y0D_lo_out[5:4],Tile_X08_Y0D_lo_out[4:3],Tile_X08_Y0D_lo_out[3:2],Tile_X08_Y0D_lo_out[2],Tile_X08_Y0D_hi_out[2:1],Tile_X08_Y0D_lo_out[0],Tile_X08_Y0D_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X08_Y0D_tile_id (
    .in(Tile_X08_Y0D_tile_id_in),
    .out(Tile_X08_Y0D_tile_id_out)
);
Tile_PE Tile_X08_Y0E (
    .SB_T0_EAST_SB_IN_B1(Tile_X09_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X09_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X08_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X08_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X08_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X08_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X08_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X08_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X08_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X08_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X08_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X08_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X07_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X07_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X08_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X08_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X09_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X09_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X08_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X08_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X08_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X08_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X08_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X08_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X08_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X08_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X08_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X08_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X07_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X07_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X08_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X08_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X09_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X09_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X08_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X08_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X08_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X08_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X08_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X08_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X08_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X08_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X08_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X08_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X07_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X07_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X08_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X08_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X09_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X09_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X08_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X08_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X08_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X08_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X08_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X08_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X08_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X08_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X08_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X08_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X07_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X07_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X08_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X08_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X09_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X09_Y0E_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X08_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X08_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X08_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X08_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X08_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X08_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X08_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X08_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X08_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X08_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X07_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X07_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X08_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X08_Y0E_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X08_Y0D_clk_out),
    .clk_out(Tile_X08_Y0E_clk_out),
    .clk_pass_through(Tile_X08_Y0D_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X08_Y0E_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X08_Y0E_clk_pass_through_out_right),
    .config_config_addr(Tile_X08_Y0D_config_out_config_addr),
    .config_config_data(Tile_X08_Y0D_config_out_config_data),
    .config_out_config_addr(Tile_X08_Y0E_config_out_config_addr),
    .config_out_config_data(Tile_X08_Y0E_config_out_config_data),
    .config_out_read(Tile_X08_Y0E_config_out_read),
    .config_out_write(Tile_X08_Y0E_config_out_write),
    .config_read(Tile_X08_Y0D_config_out_read),
    .config_write(Tile_X08_Y0D_config_out_write),
    .hi(Tile_X08_Y0E_hi_unq1),
    .lo(Tile_X08_Y0E_lo_unq1),
    .read_config_data(Tile_X08_Y0E_read_config_data),
    .read_config_data_in(Tile_X08_Y0D_read_config_data),
    .reset(Tile_X08_Y0D_reset_out),
    .reset_out(Tile_X08_Y0E_reset_out),
    .stall(Tile_X08_Y0D_stall_out),
    .stall_out(Tile_X08_Y0E_stall_out),
    .tile_id(Tile_X08_Y0E_tile_id_in)
);
mantle_wire__typeBit9 Tile_X08_Y0E_hi (
    .in(Tile_X08_Y0E_hi_unq1),
    .out(Tile_X08_Y0E_hi_out)
);
mantle_wire__typeBit8 Tile_X08_Y0E_lo (
    .in(Tile_X08_Y0E_lo_unq1),
    .out(Tile_X08_Y0E_lo_out)
);
wire [15:0] Tile_X08_Y0E_tile_id_out;
assign Tile_X08_Y0E_tile_id_out = {Tile_X08_Y0E_lo_out[7],Tile_X08_Y0E_lo_out[7:6],Tile_X08_Y0E_lo_out[6],Tile_X08_Y0E_hi_out[6],Tile_X08_Y0E_lo_out[5:4],Tile_X08_Y0E_lo_out[4:3],Tile_X08_Y0E_lo_out[3:2],Tile_X08_Y0E_lo_out[2],Tile_X08_Y0E_hi_out[2:1],Tile_X08_Y0E_hi_out[1],Tile_X08_Y0E_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X08_Y0E_tile_id (
    .in(Tile_X08_Y0E_tile_id_in),
    .out(Tile_X08_Y0E_tile_id_out)
);
Tile_PE Tile_X08_Y0F (
    .SB_T0_EAST_SB_IN_B1(Tile_X09_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X09_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X08_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X08_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X08_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X08_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X08_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X08_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X08_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X08_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X08_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X08_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X07_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X07_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X08_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X08_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X09_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X09_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X08_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X08_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X08_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X08_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X08_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X08_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X08_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X08_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X08_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X08_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X07_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X07_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X08_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X08_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X09_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X09_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X08_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X08_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X08_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X08_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X08_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X08_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X08_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X08_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X08_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X08_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X07_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X07_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X08_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X08_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X09_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X09_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X08_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X08_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X08_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X08_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X08_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X08_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X08_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X08_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X08_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X08_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X07_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X07_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X08_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X08_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X09_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X09_Y0F_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X08_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X08_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X08_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X08_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X08_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X08_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X08_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X08_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X08_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X08_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X07_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X07_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X08_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X08_Y0F_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X08_Y0E_clk_out),
    .clk_out(Tile_X08_Y0F_clk_out),
    .clk_pass_through(Tile_X08_Y0E_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X08_Y0F_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X08_Y0F_clk_pass_through_out_right),
    .config_config_addr(Tile_X08_Y0E_config_out_config_addr),
    .config_config_data(Tile_X08_Y0E_config_out_config_data),
    .config_out_config_addr(Tile_X08_Y0F_config_out_config_addr),
    .config_out_config_data(Tile_X08_Y0F_config_out_config_data),
    .config_out_read(Tile_X08_Y0F_config_out_read),
    .config_out_write(Tile_X08_Y0F_config_out_write),
    .config_read(Tile_X08_Y0E_config_out_read),
    .config_write(Tile_X08_Y0E_config_out_write),
    .hi(Tile_X08_Y0F_hi_unq1),
    .lo(Tile_X08_Y0F_lo_unq1),
    .read_config_data(Tile_X08_Y0F_read_config_data),
    .read_config_data_in(Tile_X08_Y0E_read_config_data),
    .reset(Tile_X08_Y0E_reset_out),
    .reset_out(Tile_X08_Y0F_reset_out),
    .stall(Tile_X08_Y0E_stall_out),
    .stall_out(Tile_X08_Y0F_stall_out),
    .tile_id(Tile_X08_Y0F_tile_id_in)
);
mantle_wire__typeBit9 Tile_X08_Y0F_hi (
    .in(Tile_X08_Y0F_hi_unq1),
    .out(Tile_X08_Y0F_hi_out)
);
mantle_wire__typeBit8 Tile_X08_Y0F_lo (
    .in(Tile_X08_Y0F_lo_unq1),
    .out(Tile_X08_Y0F_lo_out)
);
wire [15:0] Tile_X08_Y0F_tile_id_out;
assign Tile_X08_Y0F_tile_id_out = {Tile_X08_Y0F_lo_out[7],Tile_X08_Y0F_lo_out[7:6],Tile_X08_Y0F_lo_out[6],Tile_X08_Y0F_hi_out[6],Tile_X08_Y0F_lo_out[5:4],Tile_X08_Y0F_lo_out[4:3],Tile_X08_Y0F_lo_out[3:2],Tile_X08_Y0F_lo_out[2],Tile_X08_Y0F_hi_out[2:1],Tile_X08_Y0F_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X08_Y0F_tile_id (
    .in(Tile_X08_Y0F_tile_id_in),
    .out(Tile_X08_Y0F_tile_id_out)
);
Tile_PE Tile_X08_Y10 (
    .SB_T0_EAST_SB_IN_B1(Tile_X09_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X09_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X08_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X08_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X08_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X08_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X08_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X08_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T0_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X08_Y10_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X08_Y10_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X07_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X07_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X08_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X08_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X09_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X09_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X08_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X08_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X08_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X08_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X08_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X08_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T1_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X08_Y10_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X08_Y10_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X07_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X07_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X08_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X08_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X09_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X09_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X08_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X08_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X08_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X08_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X08_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X08_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T2_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X08_Y10_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X08_Y10_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X07_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X07_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X08_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X08_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X09_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X09_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X08_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X08_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X08_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X08_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X08_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X08_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T3_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X08_Y10_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X08_Y10_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X07_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X07_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X08_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X08_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X09_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X09_Y10_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X08_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X08_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X08_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X08_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X08_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X08_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T4_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X08_Y10_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X08_Y10_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X07_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X07_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X08_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X08_Y10_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X08_Y0F_clk_out),
    .clk_out(Tile_X08_Y10_clk_out),
    .clk_pass_through(Tile_X08_Y0F_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X08_Y10_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X08_Y10_clk_pass_through_out_right),
    .config_config_addr(Tile_X08_Y0F_config_out_config_addr),
    .config_config_data(Tile_X08_Y0F_config_out_config_data),
    .config_out_config_addr(Tile_X08_Y10_config_out_config_addr),
    .config_out_config_data(Tile_X08_Y10_config_out_config_data),
    .config_out_read(Tile_X08_Y10_config_out_read),
    .config_out_write(Tile_X08_Y10_config_out_write),
    .config_read(Tile_X08_Y0F_config_out_read),
    .config_write(Tile_X08_Y0F_config_out_write),
    .hi(Tile_X08_Y10_hi),
    .lo(Tile_X08_Y10_lo_unq1),
    .read_config_data(Tile_X08_Y10_read_config_data),
    .read_config_data_in(Tile_X08_Y0F_read_config_data),
    .reset(Tile_X08_Y0F_reset_out),
    .reset_out(Tile_X08_Y10_reset_out),
    .stall(Tile_X08_Y0F_stall_out),
    .stall_out(Tile_X08_Y10_stall_out),
    .tile_id(Tile_X08_Y10_tile_id_in)
);
mantle_wire__typeBit8 Tile_X08_Y10_lo (
    .in(Tile_X08_Y10_lo_unq1),
    .out(Tile_X08_Y10_lo_out)
);
wire [15:0] Tile_X08_Y10_tile_id_out;
assign Tile_X08_Y10_tile_id_out = {Tile_X08_Y10_lo_out[7],Tile_X08_Y10_lo_out[7:6],Tile_X08_Y10_lo_out[6],Tile_X08_Y10_hi[6],Tile_X08_Y10_lo_out[5:4],Tile_X08_Y10_lo_out[4:3],Tile_X08_Y10_lo_out[3:2],Tile_X08_Y10_hi[2],Tile_X08_Y10_lo_out[1],Tile_X08_Y10_lo_out[1:0],Tile_X08_Y10_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X08_Y10_tile_id (
    .in(Tile_X08_Y10_tile_id_in),
    .out(Tile_X08_Y10_tile_id_out)
);
wire [15:0] Tile_X09_Y00_tile_id;
assign Tile_X09_Y00_tile_id = {Tile_X09_Y00_lo[7],Tile_X09_Y00_lo[7:6],Tile_X09_Y00_lo[6],Tile_X09_Y00_hi[6],Tile_X09_Y00_lo[5:4],Tile_X09_Y00_hi[4],Tile_X09_Y00_lo[3],Tile_X09_Y00_lo[3:2],Tile_X09_Y00_lo[2:1],Tile_X09_Y00_lo[1:0],Tile_X09_Y00_lo[0]};
Tile_io_core Tile_X09_Y00 (
    .tile_id(Tile_X09_Y00_tile_id),
    .glb2io_1(glb2io_1_X09_Y00),
    .f2io_1(Tile_X09_Y01_SB_T0_NORTH_SB_OUT_B1),
    .io2glb_1(Tile_X09_Y00_io2glb_1),
    .io2f_1(Tile_X09_Y00_io2f_1),
    .glb2io_16(glb2io_16_X09_Y00),
    .f2io_16(Tile_X09_Y01_SB_T0_NORTH_SB_OUT_B16),
    .io2glb_16(Tile_X09_Y00_io2glb_16),
    .io2f_16(Tile_X09_Y00_io2f_16),
    .hi(Tile_X09_Y00_hi),
    .lo(Tile_X09_Y00_lo)
);
Tile_PE Tile_X09_Y01 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0A_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0A_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X09_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X09_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X09_Y00_io2f_1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X09_Y00_io2f_16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X09_Y01_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X09_Y01_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X09_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X09_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X09_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X09_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X08_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X08_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X09_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X09_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0A_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0A_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X09_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X09_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X09_Y00_io2f_1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X09_Y00_io2f_16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X09_Y01_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X09_Y01_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X09_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X09_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X09_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X09_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X08_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X08_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X09_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X09_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0A_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0A_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X09_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X09_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X09_Y00_io2f_1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X09_Y00_io2f_16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X09_Y01_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X09_Y01_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X09_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X09_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X09_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X09_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X08_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X08_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X09_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X09_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0A_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0A_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X09_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X09_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X09_Y00_io2f_1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X09_Y00_io2f_16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X09_Y01_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X09_Y01_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X09_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X09_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X09_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X09_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X08_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X08_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X09_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X09_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0A_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0A_Y01_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X09_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X09_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X09_Y00_io2f_1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X09_Y00_io2f_16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X09_Y01_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X09_Y01_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X09_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X09_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X09_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X09_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X08_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X08_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X09_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X09_Y01_SB_T4_WEST_SB_OUT_B16),
    .clk(clk),
    .clk_out(Tile_X09_Y01_clk_out),
    .clk_pass_through(clk),
    .clk_pass_through_out_bot(Tile_X09_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X09_Y01_clk_pass_through_out_right),
    .config_config_addr(config_9_config_addr),
    .config_config_data(config_9_config_data),
    .config_out_config_addr(Tile_X09_Y01_config_out_config_addr),
    .config_out_config_data(Tile_X09_Y01_config_out_config_data),
    .config_out_read(Tile_X09_Y01_config_out_read),
    .config_out_write(Tile_X09_Y01_config_out_write),
    .config_read(config_9_read),
    .config_write(config_9_write),
    .hi(Tile_X09_Y01_hi),
    .lo(Tile_X09_Y01_lo_unq1),
    .read_config_data(Tile_X09_Y01_read_config_data),
    .read_config_data_in(const_0_32_out),
    .reset(reset),
    .reset_out(Tile_X09_Y01_reset_out),
    .stall(stall[9]),
    .stall_out(Tile_X09_Y01_stall_out),
    .tile_id(Tile_X09_Y01_tile_id_in)
);
mantle_wire__typeBit8 Tile_X09_Y01_lo (
    .in(Tile_X09_Y01_lo_unq1),
    .out(Tile_X09_Y01_lo_out)
);
wire [15:0] Tile_X09_Y01_tile_id_out;
assign Tile_X09_Y01_tile_id_out = {Tile_X09_Y01_lo_out[7],Tile_X09_Y01_lo_out[7:6],Tile_X09_Y01_lo_out[6],Tile_X09_Y01_hi[6],Tile_X09_Y01_lo_out[5:4],Tile_X09_Y01_hi[4],Tile_X09_Y01_lo_out[3],Tile_X09_Y01_lo_out[3:2],Tile_X09_Y01_lo_out[2:1],Tile_X09_Y01_lo_out[1:0],Tile_X09_Y01_hi[0]};
mantle_wire__typeBitIn16 Tile_X09_Y01_tile_id (
    .in(Tile_X09_Y01_tile_id_in),
    .out(Tile_X09_Y01_tile_id_out)
);
Tile_PE Tile_X09_Y02 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0A_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0A_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X09_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X09_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X09_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X09_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X09_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X09_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X09_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X09_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X09_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X09_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X08_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X08_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X09_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X09_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0A_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0A_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X09_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X09_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X09_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X09_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X09_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X09_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X09_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X09_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X09_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X09_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X08_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X08_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X09_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X09_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0A_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0A_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X09_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X09_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X09_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X09_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X09_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X09_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X09_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X09_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X09_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X09_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X08_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X08_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X09_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X09_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0A_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0A_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X09_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X09_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X09_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X09_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X09_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X09_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X09_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X09_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X09_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X09_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X08_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X08_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X09_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X09_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0A_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0A_Y02_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X09_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X09_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X09_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X09_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X09_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X09_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X09_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X09_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X09_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X09_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X08_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X08_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X09_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X09_Y02_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X09_Y01_clk_out),
    .clk_out(Tile_X09_Y02_clk_out),
    .clk_pass_through(Tile_X09_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X09_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X09_Y02_clk_pass_through_out_right),
    .config_config_addr(Tile_X09_Y01_config_out_config_addr),
    .config_config_data(Tile_X09_Y01_config_out_config_data),
    .config_out_config_addr(Tile_X09_Y02_config_out_config_addr),
    .config_out_config_data(Tile_X09_Y02_config_out_config_data),
    .config_out_read(Tile_X09_Y02_config_out_read),
    .config_out_write(Tile_X09_Y02_config_out_write),
    .config_read(Tile_X09_Y01_config_out_read),
    .config_write(Tile_X09_Y01_config_out_write),
    .hi(Tile_X09_Y02_hi),
    .lo(Tile_X09_Y02_lo_unq1),
    .read_config_data(Tile_X09_Y02_read_config_data),
    .read_config_data_in(Tile_X09_Y01_read_config_data),
    .reset(Tile_X09_Y01_reset_out),
    .reset_out(Tile_X09_Y02_reset_out),
    .stall(Tile_X09_Y01_stall_out),
    .stall_out(Tile_X09_Y02_stall_out),
    .tile_id(Tile_X09_Y02_tile_id_in)
);
mantle_wire__typeBit8 Tile_X09_Y02_lo (
    .in(Tile_X09_Y02_lo_unq1),
    .out(Tile_X09_Y02_lo_out)
);
wire [15:0] Tile_X09_Y02_tile_id_out;
assign Tile_X09_Y02_tile_id_out = {Tile_X09_Y02_lo_out[7],Tile_X09_Y02_lo_out[7:6],Tile_X09_Y02_lo_out[6],Tile_X09_Y02_hi[6],Tile_X09_Y02_lo_out[5:4],Tile_X09_Y02_hi[4],Tile_X09_Y02_lo_out[3],Tile_X09_Y02_lo_out[3:2],Tile_X09_Y02_lo_out[2:1],Tile_X09_Y02_lo_out[1],Tile_X09_Y02_hi[1],Tile_X09_Y02_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X09_Y02_tile_id (
    .in(Tile_X09_Y02_tile_id_in),
    .out(Tile_X09_Y02_tile_id_out)
);
Tile_PE Tile_X09_Y03 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0A_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0A_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X09_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X09_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X09_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X09_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X09_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X09_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X09_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X09_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X09_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X09_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X08_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X08_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X09_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X09_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0A_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0A_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X09_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X09_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X09_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X09_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X09_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X09_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X09_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X09_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X09_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X09_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X08_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X08_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X09_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X09_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0A_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0A_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X09_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X09_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X09_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X09_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X09_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X09_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X09_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X09_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X09_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X09_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X08_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X08_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X09_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X09_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0A_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0A_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X09_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X09_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X09_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X09_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X09_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X09_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X09_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X09_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X09_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X09_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X08_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X08_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X09_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X09_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0A_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0A_Y03_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X09_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X09_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X09_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X09_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X09_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X09_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X09_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X09_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X09_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X09_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X08_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X08_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X09_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X09_Y03_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X09_Y02_clk_out),
    .clk_out(Tile_X09_Y03_clk_out),
    .clk_pass_through(Tile_X09_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X09_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X09_Y03_clk_pass_through_out_right),
    .config_config_addr(Tile_X09_Y02_config_out_config_addr),
    .config_config_data(Tile_X09_Y02_config_out_config_data),
    .config_out_config_addr(Tile_X09_Y03_config_out_config_addr),
    .config_out_config_data(Tile_X09_Y03_config_out_config_data),
    .config_out_read(Tile_X09_Y03_config_out_read),
    .config_out_write(Tile_X09_Y03_config_out_write),
    .config_read(Tile_X09_Y02_config_out_read),
    .config_write(Tile_X09_Y02_config_out_write),
    .hi(Tile_X09_Y03_hi_unq1),
    .lo(Tile_X09_Y03_lo_unq1),
    .read_config_data(Tile_X09_Y03_read_config_data),
    .read_config_data_in(Tile_X09_Y02_read_config_data),
    .reset(Tile_X09_Y02_reset_out),
    .reset_out(Tile_X09_Y03_reset_out),
    .stall(Tile_X09_Y02_stall_out),
    .stall_out(Tile_X09_Y03_stall_out),
    .tile_id(Tile_X09_Y03_tile_id_in)
);
mantle_wire__typeBit9 Tile_X09_Y03_hi (
    .in(Tile_X09_Y03_hi_unq1),
    .out(Tile_X09_Y03_hi_out)
);
mantle_wire__typeBit8 Tile_X09_Y03_lo (
    .in(Tile_X09_Y03_lo_unq1),
    .out(Tile_X09_Y03_lo_out)
);
wire [15:0] Tile_X09_Y03_tile_id_out;
assign Tile_X09_Y03_tile_id_out = {Tile_X09_Y03_lo_out[7],Tile_X09_Y03_lo_out[7:6],Tile_X09_Y03_lo_out[6],Tile_X09_Y03_hi_out[6],Tile_X09_Y03_lo_out[5:4],Tile_X09_Y03_hi_out[4],Tile_X09_Y03_lo_out[3],Tile_X09_Y03_lo_out[3:2],Tile_X09_Y03_lo_out[2:1],Tile_X09_Y03_lo_out[1],Tile_X09_Y03_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X09_Y03_tile_id (
    .in(Tile_X09_Y03_tile_id_in),
    .out(Tile_X09_Y03_tile_id_out)
);
Tile_PE Tile_X09_Y04 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0A_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0A_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X09_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X09_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X09_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X09_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X09_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X09_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X09_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X09_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X09_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X09_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X08_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X08_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X09_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X09_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0A_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0A_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X09_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X09_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X09_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X09_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X09_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X09_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X09_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X09_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X09_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X09_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X08_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X08_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X09_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X09_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0A_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0A_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X09_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X09_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X09_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X09_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X09_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X09_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X09_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X09_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X09_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X09_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X08_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X08_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X09_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X09_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0A_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0A_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X09_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X09_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X09_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X09_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X09_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X09_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X09_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X09_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X09_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X09_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X08_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X08_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X09_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X09_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0A_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0A_Y04_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X09_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X09_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X09_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X09_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X09_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X09_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X09_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X09_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X09_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X09_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X08_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X08_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X09_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X09_Y04_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X09_Y03_clk_out),
    .clk_out(Tile_X09_Y04_clk_out),
    .clk_pass_through(Tile_X09_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X09_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X09_Y04_clk_pass_through_out_right),
    .config_config_addr(Tile_X09_Y03_config_out_config_addr),
    .config_config_data(Tile_X09_Y03_config_out_config_data),
    .config_out_config_addr(Tile_X09_Y04_config_out_config_addr),
    .config_out_config_data(Tile_X09_Y04_config_out_config_data),
    .config_out_read(Tile_X09_Y04_config_out_read),
    .config_out_write(Tile_X09_Y04_config_out_write),
    .config_read(Tile_X09_Y03_config_out_read),
    .config_write(Tile_X09_Y03_config_out_write),
    .hi(Tile_X09_Y04_hi),
    .lo(Tile_X09_Y04_lo_unq1),
    .read_config_data(Tile_X09_Y04_read_config_data),
    .read_config_data_in(Tile_X09_Y03_read_config_data),
    .reset(Tile_X09_Y03_reset_out),
    .reset_out(Tile_X09_Y04_reset_out),
    .stall(Tile_X09_Y03_stall_out),
    .stall_out(Tile_X09_Y04_stall_out),
    .tile_id(Tile_X09_Y04_tile_id_in)
);
mantle_wire__typeBit8 Tile_X09_Y04_lo (
    .in(Tile_X09_Y04_lo_unq1),
    .out(Tile_X09_Y04_lo_out)
);
wire [15:0] Tile_X09_Y04_tile_id_out;
assign Tile_X09_Y04_tile_id_out = {Tile_X09_Y04_lo_out[7],Tile_X09_Y04_lo_out[7:6],Tile_X09_Y04_lo_out[6],Tile_X09_Y04_hi[6],Tile_X09_Y04_lo_out[5:4],Tile_X09_Y04_hi[4],Tile_X09_Y04_lo_out[3],Tile_X09_Y04_lo_out[3:2],Tile_X09_Y04_lo_out[2:1],Tile_X09_Y04_hi[1],Tile_X09_Y04_lo_out[0],Tile_X09_Y04_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X09_Y04_tile_id (
    .in(Tile_X09_Y04_tile_id_in),
    .out(Tile_X09_Y04_tile_id_out)
);
Tile_PE Tile_X09_Y05 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0A_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0A_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X09_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X09_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X09_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X09_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X09_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X09_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X09_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X09_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X09_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X09_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X08_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X08_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X09_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X09_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0A_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0A_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X09_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X09_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X09_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X09_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X09_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X09_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X09_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X09_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X09_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X09_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X08_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X08_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X09_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X09_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0A_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0A_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X09_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X09_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X09_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X09_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X09_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X09_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X09_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X09_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X09_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X09_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X08_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X08_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X09_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X09_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0A_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0A_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X09_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X09_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X09_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X09_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X09_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X09_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X09_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X09_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X09_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X09_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X08_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X08_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X09_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X09_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0A_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0A_Y05_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X09_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X09_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X09_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X09_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X09_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X09_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X09_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X09_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X09_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X09_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X08_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X08_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X09_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X09_Y05_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X09_Y04_clk_out),
    .clk_out(Tile_X09_Y05_clk_out),
    .clk_pass_through(Tile_X09_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X09_Y05_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X09_Y05_clk_pass_through_out_right),
    .config_config_addr(Tile_X09_Y04_config_out_config_addr),
    .config_config_data(Tile_X09_Y04_config_out_config_data),
    .config_out_config_addr(Tile_X09_Y05_config_out_config_addr),
    .config_out_config_data(Tile_X09_Y05_config_out_config_data),
    .config_out_read(Tile_X09_Y05_config_out_read),
    .config_out_write(Tile_X09_Y05_config_out_write),
    .config_read(Tile_X09_Y04_config_out_read),
    .config_write(Tile_X09_Y04_config_out_write),
    .hi(Tile_X09_Y05_hi),
    .lo(Tile_X09_Y05_lo_unq1),
    .read_config_data(Tile_X09_Y05_read_config_data),
    .read_config_data_in(Tile_X09_Y04_read_config_data),
    .reset(Tile_X09_Y04_reset_out),
    .reset_out(Tile_X09_Y05_reset_out),
    .stall(Tile_X09_Y04_stall_out),
    .stall_out(Tile_X09_Y05_stall_out),
    .tile_id(Tile_X09_Y05_tile_id_in)
);
mantle_wire__typeBit8 Tile_X09_Y05_lo (
    .in(Tile_X09_Y05_lo_unq1),
    .out(Tile_X09_Y05_lo_out)
);
wire [15:0] Tile_X09_Y05_tile_id_out;
assign Tile_X09_Y05_tile_id_out = {Tile_X09_Y05_lo_out[7],Tile_X09_Y05_lo_out[7:6],Tile_X09_Y05_lo_out[6],Tile_X09_Y05_hi[6],Tile_X09_Y05_lo_out[5:4],Tile_X09_Y05_hi[4],Tile_X09_Y05_lo_out[3],Tile_X09_Y05_lo_out[3:2],Tile_X09_Y05_lo_out[2:1],Tile_X09_Y05_hi[1],Tile_X09_Y05_lo_out[0],Tile_X09_Y05_hi[0]};
mantle_wire__typeBitIn16 Tile_X09_Y05_tile_id (
    .in(Tile_X09_Y05_tile_id_in),
    .out(Tile_X09_Y05_tile_id_out)
);
Tile_PE Tile_X09_Y06 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0A_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0A_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X09_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X09_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X09_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X09_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X09_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X09_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X09_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X09_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X09_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X09_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X08_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X08_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X09_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X09_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0A_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0A_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X09_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X09_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X09_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X09_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X09_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X09_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X09_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X09_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X09_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X09_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X08_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X08_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X09_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X09_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0A_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0A_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X09_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X09_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X09_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X09_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X09_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X09_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X09_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X09_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X09_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X09_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X08_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X08_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X09_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X09_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0A_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0A_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X09_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X09_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X09_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X09_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X09_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X09_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X09_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X09_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X09_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X09_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X08_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X08_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X09_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X09_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0A_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0A_Y06_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X09_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X09_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X09_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X09_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X09_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X09_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X09_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X09_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X09_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X09_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X08_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X08_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X09_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X09_Y06_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X09_Y05_clk_out),
    .clk_out(Tile_X09_Y06_clk_out),
    .clk_pass_through(Tile_X09_Y05_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X09_Y06_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X09_Y06_clk_pass_through_out_right),
    .config_config_addr(Tile_X09_Y05_config_out_config_addr),
    .config_config_data(Tile_X09_Y05_config_out_config_data),
    .config_out_config_addr(Tile_X09_Y06_config_out_config_addr),
    .config_out_config_data(Tile_X09_Y06_config_out_config_data),
    .config_out_read(Tile_X09_Y06_config_out_read),
    .config_out_write(Tile_X09_Y06_config_out_write),
    .config_read(Tile_X09_Y05_config_out_read),
    .config_write(Tile_X09_Y05_config_out_write),
    .hi(Tile_X09_Y06_hi),
    .lo(Tile_X09_Y06_lo_unq1),
    .read_config_data(Tile_X09_Y06_read_config_data),
    .read_config_data_in(Tile_X09_Y05_read_config_data),
    .reset(Tile_X09_Y05_reset_out),
    .reset_out(Tile_X09_Y06_reset_out),
    .stall(Tile_X09_Y05_stall_out),
    .stall_out(Tile_X09_Y06_stall_out),
    .tile_id(Tile_X09_Y06_tile_id_in)
);
mantle_wire__typeBit8 Tile_X09_Y06_lo (
    .in(Tile_X09_Y06_lo_unq1),
    .out(Tile_X09_Y06_lo_out)
);
wire [15:0] Tile_X09_Y06_tile_id_out;
assign Tile_X09_Y06_tile_id_out = {Tile_X09_Y06_lo_out[7],Tile_X09_Y06_lo_out[7:6],Tile_X09_Y06_lo_out[6],Tile_X09_Y06_hi[6],Tile_X09_Y06_lo_out[5:4],Tile_X09_Y06_hi[4],Tile_X09_Y06_lo_out[3],Tile_X09_Y06_lo_out[3:2],Tile_X09_Y06_lo_out[2:1],Tile_X09_Y06_hi[1],Tile_X09_Y06_hi[1],Tile_X09_Y06_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X09_Y06_tile_id (
    .in(Tile_X09_Y06_tile_id_in),
    .out(Tile_X09_Y06_tile_id_out)
);
Tile_PE Tile_X09_Y07 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0A_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0A_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X09_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X09_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X09_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X09_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X09_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X09_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X09_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X09_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X09_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X09_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X08_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X08_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X09_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X09_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0A_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0A_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X09_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X09_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X09_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X09_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X09_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X09_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X09_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X09_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X09_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X09_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X08_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X08_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X09_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X09_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0A_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0A_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X09_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X09_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X09_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X09_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X09_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X09_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X09_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X09_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X09_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X09_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X08_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X08_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X09_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X09_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0A_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0A_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X09_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X09_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X09_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X09_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X09_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X09_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X09_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X09_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X09_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X09_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X08_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X08_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X09_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X09_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0A_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0A_Y07_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X09_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X09_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X09_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X09_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X09_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X09_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X09_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X09_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X09_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X09_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X08_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X08_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X09_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X09_Y07_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X09_Y06_clk_out),
    .clk_out(Tile_X09_Y07_clk_out),
    .clk_pass_through(Tile_X09_Y06_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X09_Y07_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X09_Y07_clk_pass_through_out_right),
    .config_config_addr(Tile_X09_Y06_config_out_config_addr),
    .config_config_data(Tile_X09_Y06_config_out_config_data),
    .config_out_config_addr(Tile_X09_Y07_config_out_config_addr),
    .config_out_config_data(Tile_X09_Y07_config_out_config_data),
    .config_out_read(Tile_X09_Y07_config_out_read),
    .config_out_write(Tile_X09_Y07_config_out_write),
    .config_read(Tile_X09_Y06_config_out_read),
    .config_write(Tile_X09_Y06_config_out_write),
    .hi(Tile_X09_Y07_hi_unq1),
    .lo(Tile_X09_Y07_lo_unq1),
    .read_config_data(Tile_X09_Y07_read_config_data),
    .read_config_data_in(Tile_X09_Y06_read_config_data),
    .reset(Tile_X09_Y06_reset_out),
    .reset_out(Tile_X09_Y07_reset_out),
    .stall(Tile_X09_Y06_stall_out),
    .stall_out(Tile_X09_Y07_stall_out),
    .tile_id(Tile_X09_Y07_tile_id_in)
);
mantle_wire__typeBit9 Tile_X09_Y07_hi (
    .in(Tile_X09_Y07_hi_unq1),
    .out(Tile_X09_Y07_hi_out)
);
mantle_wire__typeBit8 Tile_X09_Y07_lo (
    .in(Tile_X09_Y07_lo_unq1),
    .out(Tile_X09_Y07_lo_out)
);
wire [15:0] Tile_X09_Y07_tile_id_out;
assign Tile_X09_Y07_tile_id_out = {Tile_X09_Y07_lo_out[7],Tile_X09_Y07_lo_out[7:6],Tile_X09_Y07_lo_out[6],Tile_X09_Y07_hi_out[6],Tile_X09_Y07_lo_out[5:4],Tile_X09_Y07_hi_out[4],Tile_X09_Y07_lo_out[3],Tile_X09_Y07_lo_out[3:2],Tile_X09_Y07_lo_out[2:1],Tile_X09_Y07_hi_out[1],Tile_X09_Y07_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X09_Y07_tile_id (
    .in(Tile_X09_Y07_tile_id_in),
    .out(Tile_X09_Y07_tile_id_out)
);
Tile_PE Tile_X09_Y08 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0A_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0A_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X09_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X09_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X09_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X09_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X09_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X09_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X09_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X09_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X09_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X09_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X08_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X08_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X09_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X09_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0A_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0A_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X09_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X09_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X09_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X09_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X09_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X09_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X09_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X09_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X09_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X09_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X08_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X08_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X09_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X09_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0A_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0A_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X09_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X09_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X09_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X09_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X09_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X09_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X09_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X09_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X09_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X09_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X08_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X08_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X09_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X09_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0A_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0A_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X09_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X09_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X09_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X09_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X09_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X09_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X09_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X09_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X09_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X09_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X08_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X08_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X09_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X09_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0A_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0A_Y08_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X09_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X09_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X09_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X09_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X09_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X09_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X09_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X09_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X09_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X09_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X08_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X08_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X09_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X09_Y08_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X09_Y07_clk_out),
    .clk_out(Tile_X09_Y08_clk_out),
    .clk_pass_through(Tile_X09_Y07_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X09_Y08_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X09_Y08_clk_pass_through_out_right),
    .config_config_addr(Tile_X09_Y07_config_out_config_addr),
    .config_config_data(Tile_X09_Y07_config_out_config_data),
    .config_out_config_addr(Tile_X09_Y08_config_out_config_addr),
    .config_out_config_data(Tile_X09_Y08_config_out_config_data),
    .config_out_read(Tile_X09_Y08_config_out_read),
    .config_out_write(Tile_X09_Y08_config_out_write),
    .config_read(Tile_X09_Y07_config_out_read),
    .config_write(Tile_X09_Y07_config_out_write),
    .hi(Tile_X09_Y08_hi),
    .lo(Tile_X09_Y08_lo_unq1),
    .read_config_data(Tile_X09_Y08_read_config_data),
    .read_config_data_in(Tile_X09_Y07_read_config_data),
    .reset(Tile_X09_Y07_reset_out),
    .reset_out(Tile_X09_Y08_reset_out),
    .stall(Tile_X09_Y07_stall_out),
    .stall_out(Tile_X09_Y08_stall_out),
    .tile_id(Tile_X09_Y08_tile_id_in)
);
mantle_wire__typeBit8 Tile_X09_Y08_lo (
    .in(Tile_X09_Y08_lo_unq1),
    .out(Tile_X09_Y08_lo_out)
);
wire [15:0] Tile_X09_Y08_tile_id_out;
assign Tile_X09_Y08_tile_id_out = {Tile_X09_Y08_lo_out[7],Tile_X09_Y08_lo_out[7:6],Tile_X09_Y08_lo_out[6],Tile_X09_Y08_hi[6],Tile_X09_Y08_lo_out[5:4],Tile_X09_Y08_hi[4],Tile_X09_Y08_lo_out[3],Tile_X09_Y08_lo_out[3:2],Tile_X09_Y08_lo_out[2],Tile_X09_Y08_hi[2],Tile_X09_Y08_lo_out[1:0],Tile_X09_Y08_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X09_Y08_tile_id (
    .in(Tile_X09_Y08_tile_id_in),
    .out(Tile_X09_Y08_tile_id_out)
);
Tile_PE Tile_X09_Y09 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0A_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0A_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X09_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X09_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X09_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X09_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X09_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X09_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X09_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X09_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X09_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X09_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X08_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X08_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X09_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X09_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0A_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0A_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X09_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X09_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X09_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X09_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X09_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X09_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X09_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X09_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X09_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X09_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X08_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X08_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X09_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X09_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0A_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0A_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X09_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X09_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X09_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X09_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X09_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X09_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X09_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X09_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X09_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X09_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X08_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X08_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X09_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X09_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0A_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0A_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X09_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X09_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X09_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X09_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X09_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X09_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X09_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X09_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X09_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X09_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X08_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X08_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X09_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X09_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0A_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0A_Y09_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X09_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X09_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X09_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X09_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X09_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X09_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X09_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X09_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X09_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X09_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X08_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X08_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X09_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X09_Y09_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X09_Y08_clk_out),
    .clk_out(Tile_X09_Y09_clk_out),
    .clk_pass_through(Tile_X09_Y08_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X09_Y09_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X09_Y09_clk_pass_through_out_right),
    .config_config_addr(ConfigPipeStage_inst9_config_out_config_addr),
    .config_config_data(ConfigPipeStage_inst9_config_out_config_data),
    .config_out_config_addr(Tile_X09_Y09_config_out_config_addr),
    .config_out_config_data(Tile_X09_Y09_config_out_config_data),
    .config_out_read(Tile_X09_Y09_config_out_read),
    .config_out_write(Tile_X09_Y09_config_out_write),
    .config_read(ConfigPipeStage_inst9_config_out_read),
    .config_write(ConfigPipeStage_inst9_config_out_write),
    .hi(Tile_X09_Y09_hi),
    .lo(Tile_X09_Y09_lo_unq1),
    .read_config_data(Tile_X09_Y09_read_config_data),
    .read_config_data_in(Tile_X09_Y08_read_config_data),
    .reset(Tile_X09_Y08_reset_out),
    .reset_out(Tile_X09_Y09_reset_out),
    .stall(Tile_X09_Y08_stall_out),
    .stall_out(Tile_X09_Y09_stall_out),
    .tile_id(Tile_X09_Y09_tile_id_in)
);
mantle_wire__typeBit8 Tile_X09_Y09_lo (
    .in(Tile_X09_Y09_lo_unq1),
    .out(Tile_X09_Y09_lo_out)
);
wire [15:0] Tile_X09_Y09_tile_id_out;
assign Tile_X09_Y09_tile_id_out = {Tile_X09_Y09_lo_out[7],Tile_X09_Y09_lo_out[7:6],Tile_X09_Y09_lo_out[6],Tile_X09_Y09_hi[6],Tile_X09_Y09_lo_out[5:4],Tile_X09_Y09_hi[4],Tile_X09_Y09_lo_out[3],Tile_X09_Y09_lo_out[3:2],Tile_X09_Y09_lo_out[2],Tile_X09_Y09_hi[2],Tile_X09_Y09_lo_out[1:0],Tile_X09_Y09_hi[0]};
mantle_wire__typeBitIn16 Tile_X09_Y09_tile_id (
    .in(Tile_X09_Y09_tile_id_in),
    .out(Tile_X09_Y09_tile_id_out)
);
Tile_PE Tile_X09_Y0A (
    .SB_T0_EAST_SB_IN_B1(Tile_X0A_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0A_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X09_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X09_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X09_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X09_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X09_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X09_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X09_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X09_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X09_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X09_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X08_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X08_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X09_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X09_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0A_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0A_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X09_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X09_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X09_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X09_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X09_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X09_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X09_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X09_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X09_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X09_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X08_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X08_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X09_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X09_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0A_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0A_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X09_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X09_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X09_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X09_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X09_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X09_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X09_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X09_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X09_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X09_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X08_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X08_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X09_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X09_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0A_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0A_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X09_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X09_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X09_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X09_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X09_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X09_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X09_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X09_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X09_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X09_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X08_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X08_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X09_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X09_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0A_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0A_Y0A_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X09_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X09_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X09_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X09_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X09_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X09_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X09_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X09_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X09_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X09_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X08_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X08_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X09_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X09_Y0A_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X09_Y09_clk_out),
    .clk_out(Tile_X09_Y0A_clk_out),
    .clk_pass_through(Tile_X09_Y09_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X09_Y0A_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X09_Y0A_clk_pass_through_out_right),
    .config_config_addr(Tile_X09_Y09_config_out_config_addr),
    .config_config_data(Tile_X09_Y09_config_out_config_data),
    .config_out_config_addr(Tile_X09_Y0A_config_out_config_addr),
    .config_out_config_data(Tile_X09_Y0A_config_out_config_data),
    .config_out_read(Tile_X09_Y0A_config_out_read),
    .config_out_write(Tile_X09_Y0A_config_out_write),
    .config_read(Tile_X09_Y09_config_out_read),
    .config_write(Tile_X09_Y09_config_out_write),
    .hi(Tile_X09_Y0A_hi),
    .lo(Tile_X09_Y0A_lo_unq1),
    .read_config_data(Tile_X09_Y0A_read_config_data),
    .read_config_data_in(Tile_X09_Y09_read_config_data),
    .reset(Tile_X09_Y09_reset_out),
    .reset_out(Tile_X09_Y0A_reset_out),
    .stall(Tile_X09_Y09_stall_out),
    .stall_out(Tile_X09_Y0A_stall_out),
    .tile_id(Tile_X09_Y0A_tile_id_in)
);
mantle_wire__typeBit8 Tile_X09_Y0A_lo (
    .in(Tile_X09_Y0A_lo_unq1),
    .out(Tile_X09_Y0A_lo_out)
);
wire [15:0] Tile_X09_Y0A_tile_id_out;
assign Tile_X09_Y0A_tile_id_out = {Tile_X09_Y0A_lo_out[7],Tile_X09_Y0A_lo_out[7:6],Tile_X09_Y0A_lo_out[6],Tile_X09_Y0A_hi[6],Tile_X09_Y0A_lo_out[5:4],Tile_X09_Y0A_hi[4],Tile_X09_Y0A_lo_out[3],Tile_X09_Y0A_lo_out[3:2],Tile_X09_Y0A_lo_out[2],Tile_X09_Y0A_hi[2],Tile_X09_Y0A_lo_out[1],Tile_X09_Y0A_hi[1],Tile_X09_Y0A_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X09_Y0A_tile_id (
    .in(Tile_X09_Y0A_tile_id_in),
    .out(Tile_X09_Y0A_tile_id_out)
);
Tile_PE Tile_X09_Y0B (
    .SB_T0_EAST_SB_IN_B1(Tile_X0A_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0A_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X09_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X09_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X09_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X09_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X09_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X09_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X09_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X09_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X09_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X09_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X08_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X08_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X09_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X09_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0A_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0A_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X09_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X09_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X09_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X09_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X09_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X09_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X09_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X09_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X09_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X09_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X08_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X08_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X09_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X09_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0A_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0A_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X09_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X09_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X09_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X09_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X09_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X09_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X09_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X09_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X09_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X09_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X08_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X08_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X09_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X09_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0A_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0A_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X09_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X09_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X09_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X09_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X09_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X09_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X09_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X09_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X09_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X09_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X08_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X08_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X09_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X09_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0A_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0A_Y0B_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X09_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X09_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X09_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X09_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X09_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X09_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X09_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X09_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X09_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X09_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X08_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X08_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X09_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X09_Y0B_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X09_Y0A_clk_out),
    .clk_out(Tile_X09_Y0B_clk_out),
    .clk_pass_through(Tile_X09_Y0A_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X09_Y0B_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X09_Y0B_clk_pass_through_out_right),
    .config_config_addr(Tile_X09_Y0A_config_out_config_addr),
    .config_config_data(Tile_X09_Y0A_config_out_config_data),
    .config_out_config_addr(Tile_X09_Y0B_config_out_config_addr),
    .config_out_config_data(Tile_X09_Y0B_config_out_config_data),
    .config_out_read(Tile_X09_Y0B_config_out_read),
    .config_out_write(Tile_X09_Y0B_config_out_write),
    .config_read(Tile_X09_Y0A_config_out_read),
    .config_write(Tile_X09_Y0A_config_out_write),
    .hi(Tile_X09_Y0B_hi_unq1),
    .lo(Tile_X09_Y0B_lo_unq1),
    .read_config_data(Tile_X09_Y0B_read_config_data),
    .read_config_data_in(Tile_X09_Y0A_read_config_data),
    .reset(Tile_X09_Y0A_reset_out),
    .reset_out(Tile_X09_Y0B_reset_out),
    .stall(Tile_X09_Y0A_stall_out),
    .stall_out(Tile_X09_Y0B_stall_out),
    .tile_id(Tile_X09_Y0B_tile_id_in)
);
mantle_wire__typeBit9 Tile_X09_Y0B_hi (
    .in(Tile_X09_Y0B_hi_unq1),
    .out(Tile_X09_Y0B_hi_out)
);
mantle_wire__typeBit8 Tile_X09_Y0B_lo (
    .in(Tile_X09_Y0B_lo_unq1),
    .out(Tile_X09_Y0B_lo_out)
);
wire [15:0] Tile_X09_Y0B_tile_id_out;
assign Tile_X09_Y0B_tile_id_out = {Tile_X09_Y0B_lo_out[7],Tile_X09_Y0B_lo_out[7:6],Tile_X09_Y0B_lo_out[6],Tile_X09_Y0B_hi_out[6],Tile_X09_Y0B_lo_out[5:4],Tile_X09_Y0B_hi_out[4],Tile_X09_Y0B_lo_out[3],Tile_X09_Y0B_lo_out[3:2],Tile_X09_Y0B_lo_out[2],Tile_X09_Y0B_hi_out[2],Tile_X09_Y0B_lo_out[1],Tile_X09_Y0B_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X09_Y0B_tile_id (
    .in(Tile_X09_Y0B_tile_id_in),
    .out(Tile_X09_Y0B_tile_id_out)
);
Tile_PE Tile_X09_Y0C (
    .SB_T0_EAST_SB_IN_B1(Tile_X0A_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0A_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X09_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X09_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X09_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X09_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X09_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X09_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X09_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X09_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X09_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X09_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X08_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X08_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X09_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X09_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0A_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0A_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X09_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X09_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X09_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X09_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X09_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X09_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X09_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X09_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X09_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X09_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X08_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X08_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X09_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X09_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0A_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0A_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X09_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X09_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X09_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X09_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X09_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X09_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X09_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X09_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X09_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X09_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X08_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X08_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X09_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X09_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0A_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0A_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X09_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X09_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X09_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X09_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X09_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X09_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X09_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X09_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X09_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X09_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X08_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X08_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X09_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X09_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0A_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0A_Y0C_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X09_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X09_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X09_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X09_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X09_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X09_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X09_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X09_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X09_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X09_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X08_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X08_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X09_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X09_Y0C_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X09_Y0B_clk_out),
    .clk_out(Tile_X09_Y0C_clk_out),
    .clk_pass_through(Tile_X09_Y0B_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X09_Y0C_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X09_Y0C_clk_pass_through_out_right),
    .config_config_addr(Tile_X09_Y0B_config_out_config_addr),
    .config_config_data(Tile_X09_Y0B_config_out_config_data),
    .config_out_config_addr(Tile_X09_Y0C_config_out_config_addr),
    .config_out_config_data(Tile_X09_Y0C_config_out_config_data),
    .config_out_read(Tile_X09_Y0C_config_out_read),
    .config_out_write(Tile_X09_Y0C_config_out_write),
    .config_read(Tile_X09_Y0B_config_out_read),
    .config_write(Tile_X09_Y0B_config_out_write),
    .hi(Tile_X09_Y0C_hi_unq1),
    .lo(Tile_X09_Y0C_lo_unq1),
    .read_config_data(Tile_X09_Y0C_read_config_data),
    .read_config_data_in(Tile_X09_Y0B_read_config_data),
    .reset(Tile_X09_Y0B_reset_out),
    .reset_out(Tile_X09_Y0C_reset_out),
    .stall(Tile_X09_Y0B_stall_out),
    .stall_out(Tile_X09_Y0C_stall_out),
    .tile_id(Tile_X09_Y0C_tile_id_in)
);
mantle_wire__typeBit9 Tile_X09_Y0C_hi (
    .in(Tile_X09_Y0C_hi_unq1),
    .out(Tile_X09_Y0C_hi_out)
);
mantle_wire__typeBit8 Tile_X09_Y0C_lo (
    .in(Tile_X09_Y0C_lo_unq1),
    .out(Tile_X09_Y0C_lo_out)
);
wire [15:0] Tile_X09_Y0C_tile_id_out;
assign Tile_X09_Y0C_tile_id_out = {Tile_X09_Y0C_lo_out[7],Tile_X09_Y0C_lo_out[7:6],Tile_X09_Y0C_lo_out[6],Tile_X09_Y0C_hi_out[6],Tile_X09_Y0C_lo_out[5:4],Tile_X09_Y0C_hi_out[4],Tile_X09_Y0C_lo_out[3],Tile_X09_Y0C_lo_out[3:2],Tile_X09_Y0C_lo_out[2],Tile_X09_Y0C_hi_out[2:1],Tile_X09_Y0C_lo_out[0],Tile_X09_Y0C_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X09_Y0C_tile_id (
    .in(Tile_X09_Y0C_tile_id_in),
    .out(Tile_X09_Y0C_tile_id_out)
);
Tile_PE Tile_X09_Y0D (
    .SB_T0_EAST_SB_IN_B1(Tile_X0A_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0A_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X09_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X09_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X09_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X09_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X09_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X09_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X09_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X09_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X09_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X09_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X08_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X08_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X09_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X09_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0A_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0A_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X09_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X09_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X09_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X09_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X09_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X09_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X09_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X09_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X09_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X09_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X08_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X08_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X09_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X09_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0A_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0A_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X09_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X09_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X09_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X09_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X09_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X09_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X09_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X09_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X09_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X09_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X08_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X08_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X09_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X09_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0A_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0A_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X09_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X09_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X09_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X09_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X09_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X09_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X09_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X09_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X09_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X09_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X08_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X08_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X09_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X09_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0A_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0A_Y0D_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X09_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X09_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X09_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X09_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X09_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X09_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X09_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X09_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X09_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X09_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X08_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X08_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X09_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X09_Y0D_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X09_Y0C_clk_out),
    .clk_out(Tile_X09_Y0D_clk_out),
    .clk_pass_through(Tile_X09_Y0C_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X09_Y0D_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X09_Y0D_clk_pass_through_out_right),
    .config_config_addr(Tile_X09_Y0C_config_out_config_addr),
    .config_config_data(Tile_X09_Y0C_config_out_config_data),
    .config_out_config_addr(Tile_X09_Y0D_config_out_config_addr),
    .config_out_config_data(Tile_X09_Y0D_config_out_config_data),
    .config_out_read(Tile_X09_Y0D_config_out_read),
    .config_out_write(Tile_X09_Y0D_config_out_write),
    .config_read(Tile_X09_Y0C_config_out_read),
    .config_write(Tile_X09_Y0C_config_out_write),
    .hi(Tile_X09_Y0D_hi_unq1),
    .lo(Tile_X09_Y0D_lo_unq1),
    .read_config_data(Tile_X09_Y0D_read_config_data),
    .read_config_data_in(Tile_X09_Y0C_read_config_data),
    .reset(Tile_X09_Y0C_reset_out),
    .reset_out(Tile_X09_Y0D_reset_out),
    .stall(Tile_X09_Y0C_stall_out),
    .stall_out(Tile_X09_Y0D_stall_out),
    .tile_id(Tile_X09_Y0D_tile_id_in)
);
mantle_wire__typeBit9 Tile_X09_Y0D_hi (
    .in(Tile_X09_Y0D_hi_unq1),
    .out(Tile_X09_Y0D_hi_out)
);
mantle_wire__typeBit8 Tile_X09_Y0D_lo (
    .in(Tile_X09_Y0D_lo_unq1),
    .out(Tile_X09_Y0D_lo_out)
);
wire [15:0] Tile_X09_Y0D_tile_id_out;
assign Tile_X09_Y0D_tile_id_out = {Tile_X09_Y0D_lo_out[7],Tile_X09_Y0D_lo_out[7:6],Tile_X09_Y0D_lo_out[6],Tile_X09_Y0D_hi_out[6],Tile_X09_Y0D_lo_out[5:4],Tile_X09_Y0D_hi_out[4],Tile_X09_Y0D_lo_out[3],Tile_X09_Y0D_lo_out[3:2],Tile_X09_Y0D_lo_out[2],Tile_X09_Y0D_hi_out[2:1],Tile_X09_Y0D_lo_out[0],Tile_X09_Y0D_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X09_Y0D_tile_id (
    .in(Tile_X09_Y0D_tile_id_in),
    .out(Tile_X09_Y0D_tile_id_out)
);
Tile_PE Tile_X09_Y0E (
    .SB_T0_EAST_SB_IN_B1(Tile_X0A_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0A_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X09_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X09_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X09_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X09_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X09_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X09_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X09_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X09_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X09_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X09_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X08_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X08_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X09_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X09_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0A_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0A_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X09_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X09_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X09_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X09_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X09_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X09_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X09_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X09_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X09_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X09_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X08_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X08_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X09_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X09_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0A_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0A_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X09_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X09_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X09_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X09_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X09_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X09_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X09_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X09_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X09_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X09_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X08_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X08_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X09_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X09_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0A_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0A_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X09_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X09_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X09_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X09_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X09_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X09_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X09_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X09_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X09_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X09_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X08_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X08_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X09_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X09_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0A_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0A_Y0E_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X09_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X09_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X09_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X09_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X09_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X09_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X09_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X09_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X09_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X09_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X08_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X08_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X09_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X09_Y0E_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X09_Y0D_clk_out),
    .clk_out(Tile_X09_Y0E_clk_out),
    .clk_pass_through(Tile_X09_Y0D_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X09_Y0E_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X09_Y0E_clk_pass_through_out_right),
    .config_config_addr(Tile_X09_Y0D_config_out_config_addr),
    .config_config_data(Tile_X09_Y0D_config_out_config_data),
    .config_out_config_addr(Tile_X09_Y0E_config_out_config_addr),
    .config_out_config_data(Tile_X09_Y0E_config_out_config_data),
    .config_out_read(Tile_X09_Y0E_config_out_read),
    .config_out_write(Tile_X09_Y0E_config_out_write),
    .config_read(Tile_X09_Y0D_config_out_read),
    .config_write(Tile_X09_Y0D_config_out_write),
    .hi(Tile_X09_Y0E_hi_unq1),
    .lo(Tile_X09_Y0E_lo_unq1),
    .read_config_data(Tile_X09_Y0E_read_config_data),
    .read_config_data_in(Tile_X09_Y0D_read_config_data),
    .reset(Tile_X09_Y0D_reset_out),
    .reset_out(Tile_X09_Y0E_reset_out),
    .stall(Tile_X09_Y0D_stall_out),
    .stall_out(Tile_X09_Y0E_stall_out),
    .tile_id(Tile_X09_Y0E_tile_id_in)
);
mantle_wire__typeBit9 Tile_X09_Y0E_hi (
    .in(Tile_X09_Y0E_hi_unq1),
    .out(Tile_X09_Y0E_hi_out)
);
mantle_wire__typeBit8 Tile_X09_Y0E_lo (
    .in(Tile_X09_Y0E_lo_unq1),
    .out(Tile_X09_Y0E_lo_out)
);
wire [15:0] Tile_X09_Y0E_tile_id_out;
assign Tile_X09_Y0E_tile_id_out = {Tile_X09_Y0E_lo_out[7],Tile_X09_Y0E_lo_out[7:6],Tile_X09_Y0E_lo_out[6],Tile_X09_Y0E_hi_out[6],Tile_X09_Y0E_lo_out[5:4],Tile_X09_Y0E_hi_out[4],Tile_X09_Y0E_lo_out[3],Tile_X09_Y0E_lo_out[3:2],Tile_X09_Y0E_lo_out[2],Tile_X09_Y0E_hi_out[2:1],Tile_X09_Y0E_hi_out[1],Tile_X09_Y0E_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X09_Y0E_tile_id (
    .in(Tile_X09_Y0E_tile_id_in),
    .out(Tile_X09_Y0E_tile_id_out)
);
Tile_PE Tile_X09_Y0F (
    .SB_T0_EAST_SB_IN_B1(Tile_X0A_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0A_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X09_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X09_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X09_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X09_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X09_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X09_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X09_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X09_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X09_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X09_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X08_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X08_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X09_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X09_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0A_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0A_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X09_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X09_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X09_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X09_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X09_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X09_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X09_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X09_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X09_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X09_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X08_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X08_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X09_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X09_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0A_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0A_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X09_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X09_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X09_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X09_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X09_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X09_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X09_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X09_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X09_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X09_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X08_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X08_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X09_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X09_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0A_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0A_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X09_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X09_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X09_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X09_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X09_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X09_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X09_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X09_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X09_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X09_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X08_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X08_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X09_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X09_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0A_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0A_Y0F_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X09_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X09_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X09_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X09_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X09_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X09_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X09_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X09_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X09_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X09_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X08_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X08_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X09_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X09_Y0F_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X09_Y0E_clk_out),
    .clk_out(Tile_X09_Y0F_clk_out),
    .clk_pass_through(Tile_X09_Y0E_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X09_Y0F_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X09_Y0F_clk_pass_through_out_right),
    .config_config_addr(Tile_X09_Y0E_config_out_config_addr),
    .config_config_data(Tile_X09_Y0E_config_out_config_data),
    .config_out_config_addr(Tile_X09_Y0F_config_out_config_addr),
    .config_out_config_data(Tile_X09_Y0F_config_out_config_data),
    .config_out_read(Tile_X09_Y0F_config_out_read),
    .config_out_write(Tile_X09_Y0F_config_out_write),
    .config_read(Tile_X09_Y0E_config_out_read),
    .config_write(Tile_X09_Y0E_config_out_write),
    .hi(Tile_X09_Y0F_hi_unq1),
    .lo(Tile_X09_Y0F_lo_unq1),
    .read_config_data(Tile_X09_Y0F_read_config_data),
    .read_config_data_in(Tile_X09_Y0E_read_config_data),
    .reset(Tile_X09_Y0E_reset_out),
    .reset_out(Tile_X09_Y0F_reset_out),
    .stall(Tile_X09_Y0E_stall_out),
    .stall_out(Tile_X09_Y0F_stall_out),
    .tile_id(Tile_X09_Y0F_tile_id_in)
);
mantle_wire__typeBit9 Tile_X09_Y0F_hi (
    .in(Tile_X09_Y0F_hi_unq1),
    .out(Tile_X09_Y0F_hi_out)
);
mantle_wire__typeBit8 Tile_X09_Y0F_lo (
    .in(Tile_X09_Y0F_lo_unq1),
    .out(Tile_X09_Y0F_lo_out)
);
wire [15:0] Tile_X09_Y0F_tile_id_out;
assign Tile_X09_Y0F_tile_id_out = {Tile_X09_Y0F_lo_out[7],Tile_X09_Y0F_lo_out[7:6],Tile_X09_Y0F_lo_out[6],Tile_X09_Y0F_hi_out[6],Tile_X09_Y0F_lo_out[5:4],Tile_X09_Y0F_hi_out[4],Tile_X09_Y0F_lo_out[3],Tile_X09_Y0F_lo_out[3:2],Tile_X09_Y0F_lo_out[2],Tile_X09_Y0F_hi_out[2:1],Tile_X09_Y0F_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X09_Y0F_tile_id (
    .in(Tile_X09_Y0F_tile_id_in),
    .out(Tile_X09_Y0F_tile_id_out)
);
Tile_PE Tile_X09_Y10 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0A_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0A_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X09_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X09_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X09_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X09_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X09_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X09_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T0_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X09_Y10_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X09_Y10_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X08_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X08_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X09_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X09_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0A_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0A_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X09_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X09_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X09_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X09_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X09_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X09_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T1_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X09_Y10_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X09_Y10_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X08_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X08_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X09_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X09_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0A_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0A_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X09_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X09_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X09_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X09_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X09_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X09_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T2_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X09_Y10_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X09_Y10_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X08_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X08_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X09_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X09_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0A_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0A_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X09_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X09_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X09_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X09_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X09_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X09_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T3_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X09_Y10_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X09_Y10_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X08_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X08_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X09_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X09_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0A_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0A_Y10_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X09_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X09_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X09_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X09_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X09_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X09_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T4_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X09_Y10_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X09_Y10_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X08_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X08_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X09_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X09_Y10_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X09_Y0F_clk_out),
    .clk_out(Tile_X09_Y10_clk_out),
    .clk_pass_through(Tile_X09_Y0F_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X09_Y10_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X09_Y10_clk_pass_through_out_right),
    .config_config_addr(Tile_X09_Y0F_config_out_config_addr),
    .config_config_data(Tile_X09_Y0F_config_out_config_data),
    .config_out_config_addr(Tile_X09_Y10_config_out_config_addr),
    .config_out_config_data(Tile_X09_Y10_config_out_config_data),
    .config_out_read(Tile_X09_Y10_config_out_read),
    .config_out_write(Tile_X09_Y10_config_out_write),
    .config_read(Tile_X09_Y0F_config_out_read),
    .config_write(Tile_X09_Y0F_config_out_write),
    .hi(Tile_X09_Y10_hi),
    .lo(Tile_X09_Y10_lo_unq1),
    .read_config_data(Tile_X09_Y10_read_config_data),
    .read_config_data_in(Tile_X09_Y0F_read_config_data),
    .reset(Tile_X09_Y0F_reset_out),
    .reset_out(Tile_X09_Y10_reset_out),
    .stall(Tile_X09_Y0F_stall_out),
    .stall_out(Tile_X09_Y10_stall_out),
    .tile_id(Tile_X09_Y10_tile_id_in)
);
mantle_wire__typeBit8 Tile_X09_Y10_lo (
    .in(Tile_X09_Y10_lo_unq1),
    .out(Tile_X09_Y10_lo_out)
);
wire [15:0] Tile_X09_Y10_tile_id_out;
assign Tile_X09_Y10_tile_id_out = {Tile_X09_Y10_lo_out[7],Tile_X09_Y10_lo_out[7:6],Tile_X09_Y10_lo_out[6],Tile_X09_Y10_hi[6],Tile_X09_Y10_lo_out[5:4],Tile_X09_Y10_hi[4],Tile_X09_Y10_lo_out[3],Tile_X09_Y10_lo_out[3:2],Tile_X09_Y10_hi[2],Tile_X09_Y10_lo_out[1],Tile_X09_Y10_lo_out[1:0],Tile_X09_Y10_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X09_Y10_tile_id (
    .in(Tile_X09_Y10_tile_id_in),
    .out(Tile_X09_Y10_tile_id_out)
);
wire [15:0] Tile_X0A_Y00_tile_id;
assign Tile_X0A_Y00_tile_id = {Tile_X0A_Y00_lo[7],Tile_X0A_Y00_lo[7:6],Tile_X0A_Y00_lo[6],Tile_X0A_Y00_hi[6],Tile_X0A_Y00_lo[5],Tile_X0A_Y00_hi[5],Tile_X0A_Y00_lo[4:3],Tile_X0A_Y00_lo[3:2],Tile_X0A_Y00_lo[2:1],Tile_X0A_Y00_lo[1:0],Tile_X0A_Y00_lo[0]};
Tile_io_core Tile_X0A_Y00 (
    .tile_id(Tile_X0A_Y00_tile_id),
    .glb2io_1(glb2io_1_X0A_Y00),
    .f2io_1(Tile_X0A_Y01_SB_T0_NORTH_SB_OUT_B1),
    .io2glb_1(Tile_X0A_Y00_io2glb_1),
    .io2f_1(Tile_X0A_Y00_io2f_1),
    .glb2io_16(glb2io_16_X0A_Y00),
    .f2io_16(Tile_X0A_Y01_SB_T0_NORTH_SB_OUT_B16),
    .io2glb_16(Tile_X0A_Y00_io2glb_16),
    .io2f_16(Tile_X0A_Y00_io2f_16),
    .hi(Tile_X0A_Y00_hi),
    .lo(Tile_X0A_Y00_lo)
);
Tile_PE Tile_X0A_Y01 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0B_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0B_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0A_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0A_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0A_Y00_io2f_1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0A_Y00_io2f_16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0A_Y01_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0A_Y01_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0A_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0A_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0A_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0A_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X09_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X09_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0A_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0A_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0B_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0B_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0A_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0A_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0A_Y00_io2f_1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0A_Y00_io2f_16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0A_Y01_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0A_Y01_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0A_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0A_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0A_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0A_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X09_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X09_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0A_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0A_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0B_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0B_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0A_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0A_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0A_Y00_io2f_1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0A_Y00_io2f_16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0A_Y01_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0A_Y01_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0A_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0A_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0A_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0A_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X09_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X09_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0A_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0A_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0B_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0B_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0A_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0A_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0A_Y00_io2f_1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0A_Y00_io2f_16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0A_Y01_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0A_Y01_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0A_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0A_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0A_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0A_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X09_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X09_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0A_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0A_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0B_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0B_Y01_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0A_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0A_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0A_Y00_io2f_1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0A_Y00_io2f_16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0A_Y01_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0A_Y01_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0A_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0A_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0A_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0A_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X09_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X09_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0A_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0A_Y01_SB_T4_WEST_SB_OUT_B16),
    .clk(clk),
    .clk_out(Tile_X0A_Y01_clk_out),
    .clk_pass_through(clk),
    .clk_pass_through_out_bot(Tile_X0A_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0A_Y01_clk_pass_through_out_right),
    .config_config_addr(config_10_config_addr),
    .config_config_data(config_10_config_data),
    .config_out_config_addr(Tile_X0A_Y01_config_out_config_addr),
    .config_out_config_data(Tile_X0A_Y01_config_out_config_data),
    .config_out_read(Tile_X0A_Y01_config_out_read),
    .config_out_write(Tile_X0A_Y01_config_out_write),
    .config_read(config_10_read),
    .config_write(config_10_write),
    .hi(Tile_X0A_Y01_hi),
    .lo(Tile_X0A_Y01_lo_unq1),
    .read_config_data(Tile_X0A_Y01_read_config_data),
    .read_config_data_in(const_0_32_out),
    .reset(reset),
    .reset_out(Tile_X0A_Y01_reset_out),
    .stall(stall[10]),
    .stall_out(Tile_X0A_Y01_stall_out),
    .tile_id(Tile_X0A_Y01_tile_id_in)
);
mantle_wire__typeBit8 Tile_X0A_Y01_lo (
    .in(Tile_X0A_Y01_lo_unq1),
    .out(Tile_X0A_Y01_lo_out)
);
wire [15:0] Tile_X0A_Y01_tile_id_out;
assign Tile_X0A_Y01_tile_id_out = {Tile_X0A_Y01_lo_out[7],Tile_X0A_Y01_lo_out[7:6],Tile_X0A_Y01_lo_out[6],Tile_X0A_Y01_hi[6],Tile_X0A_Y01_lo_out[5],Tile_X0A_Y01_hi[5],Tile_X0A_Y01_lo_out[4:3],Tile_X0A_Y01_lo_out[3:2],Tile_X0A_Y01_lo_out[2:1],Tile_X0A_Y01_lo_out[1:0],Tile_X0A_Y01_hi[0]};
mantle_wire__typeBitIn16 Tile_X0A_Y01_tile_id (
    .in(Tile_X0A_Y01_tile_id_in),
    .out(Tile_X0A_Y01_tile_id_out)
);
Tile_PE Tile_X0A_Y02 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0B_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0B_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0A_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0A_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0A_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0A_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0A_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0A_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0A_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0A_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0A_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0A_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X09_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X09_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0A_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0A_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0B_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0B_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0A_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0A_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0A_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0A_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0A_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0A_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0A_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0A_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0A_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0A_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X09_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X09_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0A_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0A_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0B_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0B_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0A_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0A_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0A_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0A_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0A_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0A_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0A_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0A_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0A_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0A_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X09_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X09_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0A_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0A_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0B_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0B_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0A_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0A_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0A_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0A_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0A_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0A_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0A_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0A_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0A_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0A_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X09_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X09_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0A_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0A_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0B_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0B_Y02_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0A_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0A_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0A_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0A_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0A_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0A_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0A_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0A_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0A_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0A_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X09_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X09_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0A_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0A_Y02_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y01_clk_out),
    .clk_out(Tile_X0A_Y02_clk_out),
    .clk_pass_through(Tile_X0A_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0A_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0A_Y02_clk_pass_through_out_right),
    .config_config_addr(Tile_X0A_Y01_config_out_config_addr),
    .config_config_data(Tile_X0A_Y01_config_out_config_data),
    .config_out_config_addr(Tile_X0A_Y02_config_out_config_addr),
    .config_out_config_data(Tile_X0A_Y02_config_out_config_data),
    .config_out_read(Tile_X0A_Y02_config_out_read),
    .config_out_write(Tile_X0A_Y02_config_out_write),
    .config_read(Tile_X0A_Y01_config_out_read),
    .config_write(Tile_X0A_Y01_config_out_write),
    .hi(Tile_X0A_Y02_hi),
    .lo(Tile_X0A_Y02_lo_unq1),
    .read_config_data(Tile_X0A_Y02_read_config_data),
    .read_config_data_in(Tile_X0A_Y01_read_config_data),
    .reset(Tile_X0A_Y01_reset_out),
    .reset_out(Tile_X0A_Y02_reset_out),
    .stall(Tile_X0A_Y01_stall_out),
    .stall_out(Tile_X0A_Y02_stall_out),
    .tile_id(Tile_X0A_Y02_tile_id_in)
);
mantle_wire__typeBit8 Tile_X0A_Y02_lo (
    .in(Tile_X0A_Y02_lo_unq1),
    .out(Tile_X0A_Y02_lo_out)
);
wire [15:0] Tile_X0A_Y02_tile_id_out;
assign Tile_X0A_Y02_tile_id_out = {Tile_X0A_Y02_lo_out[7],Tile_X0A_Y02_lo_out[7:6],Tile_X0A_Y02_lo_out[6],Tile_X0A_Y02_hi[6],Tile_X0A_Y02_lo_out[5],Tile_X0A_Y02_hi[5],Tile_X0A_Y02_lo_out[4:3],Tile_X0A_Y02_lo_out[3:2],Tile_X0A_Y02_lo_out[2:1],Tile_X0A_Y02_lo_out[1],Tile_X0A_Y02_hi[1],Tile_X0A_Y02_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0A_Y02_tile_id (
    .in(Tile_X0A_Y02_tile_id_in),
    .out(Tile_X0A_Y02_tile_id_out)
);
Tile_PE Tile_X0A_Y03 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0B_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0B_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0A_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0A_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0A_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0A_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0A_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0A_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0A_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0A_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0A_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0A_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X09_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X09_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0A_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0A_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0B_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0B_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0A_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0A_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0A_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0A_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0A_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0A_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0A_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0A_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0A_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0A_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X09_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X09_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0A_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0A_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0B_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0B_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0A_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0A_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0A_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0A_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0A_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0A_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0A_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0A_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0A_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0A_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X09_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X09_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0A_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0A_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0B_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0B_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0A_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0A_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0A_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0A_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0A_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0A_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0A_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0A_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0A_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0A_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X09_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X09_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0A_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0A_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0B_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0B_Y03_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0A_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0A_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0A_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0A_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0A_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0A_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0A_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0A_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0A_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0A_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X09_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X09_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0A_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0A_Y03_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y02_clk_out),
    .clk_out(Tile_X0A_Y03_clk_out),
    .clk_pass_through(Tile_X0A_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0A_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0A_Y03_clk_pass_through_out_right),
    .config_config_addr(Tile_X0A_Y02_config_out_config_addr),
    .config_config_data(Tile_X0A_Y02_config_out_config_data),
    .config_out_config_addr(Tile_X0A_Y03_config_out_config_addr),
    .config_out_config_data(Tile_X0A_Y03_config_out_config_data),
    .config_out_read(Tile_X0A_Y03_config_out_read),
    .config_out_write(Tile_X0A_Y03_config_out_write),
    .config_read(Tile_X0A_Y02_config_out_read),
    .config_write(Tile_X0A_Y02_config_out_write),
    .hi(Tile_X0A_Y03_hi_unq1),
    .lo(Tile_X0A_Y03_lo_unq1),
    .read_config_data(Tile_X0A_Y03_read_config_data),
    .read_config_data_in(Tile_X0A_Y02_read_config_data),
    .reset(Tile_X0A_Y02_reset_out),
    .reset_out(Tile_X0A_Y03_reset_out),
    .stall(Tile_X0A_Y02_stall_out),
    .stall_out(Tile_X0A_Y03_stall_out),
    .tile_id(Tile_X0A_Y03_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0A_Y03_hi (
    .in(Tile_X0A_Y03_hi_unq1),
    .out(Tile_X0A_Y03_hi_out)
);
mantle_wire__typeBit8 Tile_X0A_Y03_lo (
    .in(Tile_X0A_Y03_lo_unq1),
    .out(Tile_X0A_Y03_lo_out)
);
wire [15:0] Tile_X0A_Y03_tile_id_out;
assign Tile_X0A_Y03_tile_id_out = {Tile_X0A_Y03_lo_out[7],Tile_X0A_Y03_lo_out[7:6],Tile_X0A_Y03_lo_out[6],Tile_X0A_Y03_hi_out[6],Tile_X0A_Y03_lo_out[5],Tile_X0A_Y03_hi_out[5],Tile_X0A_Y03_lo_out[4:3],Tile_X0A_Y03_lo_out[3:2],Tile_X0A_Y03_lo_out[2:1],Tile_X0A_Y03_lo_out[1],Tile_X0A_Y03_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X0A_Y03_tile_id (
    .in(Tile_X0A_Y03_tile_id_in),
    .out(Tile_X0A_Y03_tile_id_out)
);
Tile_PE Tile_X0A_Y04 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0B_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0B_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0A_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0A_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0A_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0A_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0A_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0A_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0A_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0A_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0A_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0A_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X09_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X09_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0A_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0A_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0B_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0B_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0A_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0A_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0A_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0A_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0A_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0A_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0A_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0A_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0A_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0A_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X09_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X09_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0A_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0A_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0B_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0B_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0A_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0A_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0A_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0A_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0A_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0A_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0A_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0A_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0A_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0A_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X09_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X09_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0A_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0A_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0B_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0B_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0A_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0A_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0A_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0A_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0A_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0A_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0A_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0A_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0A_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0A_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X09_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X09_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0A_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0A_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0B_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0B_Y04_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0A_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0A_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0A_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0A_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0A_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0A_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0A_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0A_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0A_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0A_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X09_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X09_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0A_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0A_Y04_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y03_clk_out),
    .clk_out(Tile_X0A_Y04_clk_out),
    .clk_pass_through(Tile_X0A_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0A_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0A_Y04_clk_pass_through_out_right),
    .config_config_addr(Tile_X0A_Y03_config_out_config_addr),
    .config_config_data(Tile_X0A_Y03_config_out_config_data),
    .config_out_config_addr(Tile_X0A_Y04_config_out_config_addr),
    .config_out_config_data(Tile_X0A_Y04_config_out_config_data),
    .config_out_read(Tile_X0A_Y04_config_out_read),
    .config_out_write(Tile_X0A_Y04_config_out_write),
    .config_read(Tile_X0A_Y03_config_out_read),
    .config_write(Tile_X0A_Y03_config_out_write),
    .hi(Tile_X0A_Y04_hi),
    .lo(Tile_X0A_Y04_lo_unq1),
    .read_config_data(Tile_X0A_Y04_read_config_data),
    .read_config_data_in(Tile_X0A_Y03_read_config_data),
    .reset(Tile_X0A_Y03_reset_out),
    .reset_out(Tile_X0A_Y04_reset_out),
    .stall(Tile_X0A_Y03_stall_out),
    .stall_out(Tile_X0A_Y04_stall_out),
    .tile_id(Tile_X0A_Y04_tile_id_in)
);
mantle_wire__typeBit8 Tile_X0A_Y04_lo (
    .in(Tile_X0A_Y04_lo_unq1),
    .out(Tile_X0A_Y04_lo_out)
);
wire [15:0] Tile_X0A_Y04_tile_id_out;
assign Tile_X0A_Y04_tile_id_out = {Tile_X0A_Y04_lo_out[7],Tile_X0A_Y04_lo_out[7:6],Tile_X0A_Y04_lo_out[6],Tile_X0A_Y04_hi[6],Tile_X0A_Y04_lo_out[5],Tile_X0A_Y04_hi[5],Tile_X0A_Y04_lo_out[4:3],Tile_X0A_Y04_lo_out[3:2],Tile_X0A_Y04_lo_out[2:1],Tile_X0A_Y04_hi[1],Tile_X0A_Y04_lo_out[0],Tile_X0A_Y04_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0A_Y04_tile_id (
    .in(Tile_X0A_Y04_tile_id_in),
    .out(Tile_X0A_Y04_tile_id_out)
);
Tile_PE Tile_X0A_Y05 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0B_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0B_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0A_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0A_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0A_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0A_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0A_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0A_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0A_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0A_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0A_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0A_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X09_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X09_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0A_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0A_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0B_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0B_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0A_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0A_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0A_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0A_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0A_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0A_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0A_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0A_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0A_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0A_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X09_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X09_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0A_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0A_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0B_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0B_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0A_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0A_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0A_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0A_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0A_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0A_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0A_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0A_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0A_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0A_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X09_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X09_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0A_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0A_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0B_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0B_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0A_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0A_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0A_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0A_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0A_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0A_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0A_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0A_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0A_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0A_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X09_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X09_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0A_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0A_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0B_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0B_Y05_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0A_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0A_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0A_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0A_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0A_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0A_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0A_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0A_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0A_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0A_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X09_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X09_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0A_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0A_Y05_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y04_clk_out),
    .clk_out(Tile_X0A_Y05_clk_out),
    .clk_pass_through(Tile_X0A_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0A_Y05_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0A_Y05_clk_pass_through_out_right),
    .config_config_addr(Tile_X0A_Y04_config_out_config_addr),
    .config_config_data(Tile_X0A_Y04_config_out_config_data),
    .config_out_config_addr(Tile_X0A_Y05_config_out_config_addr),
    .config_out_config_data(Tile_X0A_Y05_config_out_config_data),
    .config_out_read(Tile_X0A_Y05_config_out_read),
    .config_out_write(Tile_X0A_Y05_config_out_write),
    .config_read(Tile_X0A_Y04_config_out_read),
    .config_write(Tile_X0A_Y04_config_out_write),
    .hi(Tile_X0A_Y05_hi),
    .lo(Tile_X0A_Y05_lo_unq1),
    .read_config_data(Tile_X0A_Y05_read_config_data),
    .read_config_data_in(Tile_X0A_Y04_read_config_data),
    .reset(Tile_X0A_Y04_reset_out),
    .reset_out(Tile_X0A_Y05_reset_out),
    .stall(Tile_X0A_Y04_stall_out),
    .stall_out(Tile_X0A_Y05_stall_out),
    .tile_id(Tile_X0A_Y05_tile_id_in)
);
mantle_wire__typeBit8 Tile_X0A_Y05_lo (
    .in(Tile_X0A_Y05_lo_unq1),
    .out(Tile_X0A_Y05_lo_out)
);
wire [15:0] Tile_X0A_Y05_tile_id_out;
assign Tile_X0A_Y05_tile_id_out = {Tile_X0A_Y05_lo_out[7],Tile_X0A_Y05_lo_out[7:6],Tile_X0A_Y05_lo_out[6],Tile_X0A_Y05_hi[6],Tile_X0A_Y05_lo_out[5],Tile_X0A_Y05_hi[5],Tile_X0A_Y05_lo_out[4:3],Tile_X0A_Y05_lo_out[3:2],Tile_X0A_Y05_lo_out[2:1],Tile_X0A_Y05_hi[1],Tile_X0A_Y05_lo_out[0],Tile_X0A_Y05_hi[0]};
mantle_wire__typeBitIn16 Tile_X0A_Y05_tile_id (
    .in(Tile_X0A_Y05_tile_id_in),
    .out(Tile_X0A_Y05_tile_id_out)
);
Tile_PE Tile_X0A_Y06 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0B_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0B_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0A_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0A_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0A_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0A_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0A_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0A_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0A_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0A_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0A_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0A_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X09_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X09_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0A_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0A_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0B_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0B_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0A_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0A_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0A_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0A_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0A_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0A_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0A_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0A_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0A_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0A_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X09_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X09_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0A_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0A_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0B_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0B_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0A_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0A_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0A_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0A_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0A_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0A_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0A_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0A_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0A_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0A_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X09_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X09_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0A_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0A_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0B_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0B_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0A_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0A_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0A_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0A_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0A_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0A_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0A_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0A_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0A_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0A_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X09_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X09_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0A_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0A_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0B_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0B_Y06_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0A_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0A_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0A_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0A_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0A_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0A_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0A_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0A_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0A_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0A_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X09_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X09_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0A_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0A_Y06_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y05_clk_out),
    .clk_out(Tile_X0A_Y06_clk_out),
    .clk_pass_through(Tile_X0A_Y05_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0A_Y06_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0A_Y06_clk_pass_through_out_right),
    .config_config_addr(Tile_X0A_Y05_config_out_config_addr),
    .config_config_data(Tile_X0A_Y05_config_out_config_data),
    .config_out_config_addr(Tile_X0A_Y06_config_out_config_addr),
    .config_out_config_data(Tile_X0A_Y06_config_out_config_data),
    .config_out_read(Tile_X0A_Y06_config_out_read),
    .config_out_write(Tile_X0A_Y06_config_out_write),
    .config_read(Tile_X0A_Y05_config_out_read),
    .config_write(Tile_X0A_Y05_config_out_write),
    .hi(Tile_X0A_Y06_hi),
    .lo(Tile_X0A_Y06_lo_unq1),
    .read_config_data(Tile_X0A_Y06_read_config_data),
    .read_config_data_in(Tile_X0A_Y05_read_config_data),
    .reset(Tile_X0A_Y05_reset_out),
    .reset_out(Tile_X0A_Y06_reset_out),
    .stall(Tile_X0A_Y05_stall_out),
    .stall_out(Tile_X0A_Y06_stall_out),
    .tile_id(Tile_X0A_Y06_tile_id_in)
);
mantle_wire__typeBit8 Tile_X0A_Y06_lo (
    .in(Tile_X0A_Y06_lo_unq1),
    .out(Tile_X0A_Y06_lo_out)
);
wire [15:0] Tile_X0A_Y06_tile_id_out;
assign Tile_X0A_Y06_tile_id_out = {Tile_X0A_Y06_lo_out[7],Tile_X0A_Y06_lo_out[7:6],Tile_X0A_Y06_lo_out[6],Tile_X0A_Y06_hi[6],Tile_X0A_Y06_lo_out[5],Tile_X0A_Y06_hi[5],Tile_X0A_Y06_lo_out[4:3],Tile_X0A_Y06_lo_out[3:2],Tile_X0A_Y06_lo_out[2:1],Tile_X0A_Y06_hi[1],Tile_X0A_Y06_hi[1],Tile_X0A_Y06_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0A_Y06_tile_id (
    .in(Tile_X0A_Y06_tile_id_in),
    .out(Tile_X0A_Y06_tile_id_out)
);
Tile_PE Tile_X0A_Y07 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0B_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0B_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0A_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0A_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0A_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0A_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0A_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0A_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0A_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0A_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0A_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0A_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X09_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X09_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0A_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0A_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0B_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0B_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0A_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0A_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0A_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0A_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0A_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0A_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0A_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0A_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0A_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0A_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X09_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X09_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0A_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0A_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0B_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0B_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0A_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0A_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0A_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0A_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0A_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0A_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0A_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0A_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0A_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0A_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X09_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X09_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0A_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0A_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0B_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0B_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0A_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0A_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0A_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0A_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0A_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0A_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0A_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0A_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0A_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0A_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X09_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X09_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0A_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0A_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0B_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0B_Y07_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0A_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0A_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0A_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0A_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0A_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0A_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0A_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0A_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0A_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0A_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X09_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X09_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0A_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0A_Y07_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y06_clk_out),
    .clk_out(Tile_X0A_Y07_clk_out),
    .clk_pass_through(Tile_X0A_Y06_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0A_Y07_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0A_Y07_clk_pass_through_out_right),
    .config_config_addr(Tile_X0A_Y06_config_out_config_addr),
    .config_config_data(Tile_X0A_Y06_config_out_config_data),
    .config_out_config_addr(Tile_X0A_Y07_config_out_config_addr),
    .config_out_config_data(Tile_X0A_Y07_config_out_config_data),
    .config_out_read(Tile_X0A_Y07_config_out_read),
    .config_out_write(Tile_X0A_Y07_config_out_write),
    .config_read(Tile_X0A_Y06_config_out_read),
    .config_write(Tile_X0A_Y06_config_out_write),
    .hi(Tile_X0A_Y07_hi_unq1),
    .lo(Tile_X0A_Y07_lo_unq1),
    .read_config_data(Tile_X0A_Y07_read_config_data),
    .read_config_data_in(Tile_X0A_Y06_read_config_data),
    .reset(Tile_X0A_Y06_reset_out),
    .reset_out(Tile_X0A_Y07_reset_out),
    .stall(Tile_X0A_Y06_stall_out),
    .stall_out(Tile_X0A_Y07_stall_out),
    .tile_id(Tile_X0A_Y07_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0A_Y07_hi (
    .in(Tile_X0A_Y07_hi_unq1),
    .out(Tile_X0A_Y07_hi_out)
);
mantle_wire__typeBit8 Tile_X0A_Y07_lo (
    .in(Tile_X0A_Y07_lo_unq1),
    .out(Tile_X0A_Y07_lo_out)
);
wire [15:0] Tile_X0A_Y07_tile_id_out;
assign Tile_X0A_Y07_tile_id_out = {Tile_X0A_Y07_lo_out[7],Tile_X0A_Y07_lo_out[7:6],Tile_X0A_Y07_lo_out[6],Tile_X0A_Y07_hi_out[6],Tile_X0A_Y07_lo_out[5],Tile_X0A_Y07_hi_out[5],Tile_X0A_Y07_lo_out[4:3],Tile_X0A_Y07_lo_out[3:2],Tile_X0A_Y07_lo_out[2:1],Tile_X0A_Y07_hi_out[1],Tile_X0A_Y07_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X0A_Y07_tile_id (
    .in(Tile_X0A_Y07_tile_id_in),
    .out(Tile_X0A_Y07_tile_id_out)
);
Tile_PE Tile_X0A_Y08 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0B_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0B_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0A_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0A_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0A_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0A_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0A_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0A_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0A_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0A_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0A_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0A_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X09_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X09_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0A_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0A_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0B_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0B_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0A_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0A_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0A_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0A_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0A_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0A_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0A_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0A_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0A_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0A_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X09_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X09_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0A_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0A_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0B_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0B_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0A_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0A_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0A_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0A_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0A_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0A_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0A_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0A_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0A_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0A_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X09_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X09_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0A_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0A_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0B_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0B_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0A_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0A_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0A_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0A_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0A_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0A_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0A_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0A_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0A_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0A_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X09_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X09_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0A_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0A_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0B_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0B_Y08_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0A_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0A_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0A_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0A_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0A_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0A_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0A_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0A_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0A_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0A_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X09_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X09_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0A_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0A_Y08_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y07_clk_out),
    .clk_out(Tile_X0A_Y08_clk_out),
    .clk_pass_through(Tile_X0A_Y07_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0A_Y08_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0A_Y08_clk_pass_through_out_right),
    .config_config_addr(Tile_X0A_Y07_config_out_config_addr),
    .config_config_data(Tile_X0A_Y07_config_out_config_data),
    .config_out_config_addr(Tile_X0A_Y08_config_out_config_addr),
    .config_out_config_data(Tile_X0A_Y08_config_out_config_data),
    .config_out_read(Tile_X0A_Y08_config_out_read),
    .config_out_write(Tile_X0A_Y08_config_out_write),
    .config_read(Tile_X0A_Y07_config_out_read),
    .config_write(Tile_X0A_Y07_config_out_write),
    .hi(Tile_X0A_Y08_hi),
    .lo(Tile_X0A_Y08_lo_unq1),
    .read_config_data(Tile_X0A_Y08_read_config_data),
    .read_config_data_in(Tile_X0A_Y07_read_config_data),
    .reset(Tile_X0A_Y07_reset_out),
    .reset_out(Tile_X0A_Y08_reset_out),
    .stall(Tile_X0A_Y07_stall_out),
    .stall_out(Tile_X0A_Y08_stall_out),
    .tile_id(Tile_X0A_Y08_tile_id_in)
);
mantle_wire__typeBit8 Tile_X0A_Y08_lo (
    .in(Tile_X0A_Y08_lo_unq1),
    .out(Tile_X0A_Y08_lo_out)
);
wire [15:0] Tile_X0A_Y08_tile_id_out;
assign Tile_X0A_Y08_tile_id_out = {Tile_X0A_Y08_lo_out[7],Tile_X0A_Y08_lo_out[7:6],Tile_X0A_Y08_lo_out[6],Tile_X0A_Y08_hi[6],Tile_X0A_Y08_lo_out[5],Tile_X0A_Y08_hi[5],Tile_X0A_Y08_lo_out[4:3],Tile_X0A_Y08_lo_out[3:2],Tile_X0A_Y08_lo_out[2],Tile_X0A_Y08_hi[2],Tile_X0A_Y08_lo_out[1:0],Tile_X0A_Y08_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0A_Y08_tile_id (
    .in(Tile_X0A_Y08_tile_id_in),
    .out(Tile_X0A_Y08_tile_id_out)
);
Tile_PE Tile_X0A_Y09 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0B_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0B_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0A_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0A_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0A_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0A_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0A_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0A_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0A_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0A_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0A_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0A_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X09_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X09_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0A_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0A_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0B_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0B_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0A_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0A_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0A_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0A_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0A_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0A_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0A_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0A_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0A_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0A_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X09_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X09_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0A_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0A_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0B_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0B_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0A_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0A_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0A_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0A_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0A_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0A_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0A_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0A_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0A_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0A_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X09_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X09_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0A_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0A_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0B_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0B_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0A_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0A_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0A_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0A_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0A_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0A_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0A_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0A_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0A_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0A_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X09_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X09_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0A_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0A_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0B_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0B_Y09_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0A_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0A_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0A_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0A_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0A_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0A_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0A_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0A_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0A_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0A_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X09_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X09_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0A_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0A_Y09_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y08_clk_out),
    .clk_out(Tile_X0A_Y09_clk_out),
    .clk_pass_through(Tile_X0A_Y08_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0A_Y09_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0A_Y09_clk_pass_through_out_right),
    .config_config_addr(ConfigPipeStage_inst10_config_out_config_addr),
    .config_config_data(ConfigPipeStage_inst10_config_out_config_data),
    .config_out_config_addr(Tile_X0A_Y09_config_out_config_addr),
    .config_out_config_data(Tile_X0A_Y09_config_out_config_data),
    .config_out_read(Tile_X0A_Y09_config_out_read),
    .config_out_write(Tile_X0A_Y09_config_out_write),
    .config_read(ConfigPipeStage_inst10_config_out_read),
    .config_write(ConfigPipeStage_inst10_config_out_write),
    .hi(Tile_X0A_Y09_hi),
    .lo(Tile_X0A_Y09_lo_unq1),
    .read_config_data(Tile_X0A_Y09_read_config_data),
    .read_config_data_in(Tile_X0A_Y08_read_config_data),
    .reset(Tile_X0A_Y08_reset_out),
    .reset_out(Tile_X0A_Y09_reset_out),
    .stall(Tile_X0A_Y08_stall_out),
    .stall_out(Tile_X0A_Y09_stall_out),
    .tile_id(Tile_X0A_Y09_tile_id_in)
);
mantle_wire__typeBit8 Tile_X0A_Y09_lo (
    .in(Tile_X0A_Y09_lo_unq1),
    .out(Tile_X0A_Y09_lo_out)
);
wire [15:0] Tile_X0A_Y09_tile_id_out;
assign Tile_X0A_Y09_tile_id_out = {Tile_X0A_Y09_lo_out[7],Tile_X0A_Y09_lo_out[7:6],Tile_X0A_Y09_lo_out[6],Tile_X0A_Y09_hi[6],Tile_X0A_Y09_lo_out[5],Tile_X0A_Y09_hi[5],Tile_X0A_Y09_lo_out[4:3],Tile_X0A_Y09_lo_out[3:2],Tile_X0A_Y09_lo_out[2],Tile_X0A_Y09_hi[2],Tile_X0A_Y09_lo_out[1:0],Tile_X0A_Y09_hi[0]};
mantle_wire__typeBitIn16 Tile_X0A_Y09_tile_id (
    .in(Tile_X0A_Y09_tile_id_in),
    .out(Tile_X0A_Y09_tile_id_out)
);
Tile_PE Tile_X0A_Y0A (
    .SB_T0_EAST_SB_IN_B1(Tile_X0B_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0B_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0A_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0A_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0A_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0A_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0A_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0A_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0A_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0A_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0A_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0A_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X09_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X09_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0A_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0A_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0B_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0B_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0A_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0A_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0A_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0A_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0A_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0A_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0A_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0A_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0A_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0A_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X09_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X09_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0A_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0A_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0B_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0B_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0A_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0A_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0A_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0A_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0A_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0A_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0A_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0A_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0A_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0A_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X09_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X09_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0A_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0A_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0B_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0B_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0A_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0A_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0A_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0A_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0A_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0A_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0A_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0A_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0A_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0A_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X09_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X09_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0A_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0A_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0B_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0B_Y0A_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0A_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0A_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0A_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0A_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0A_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0A_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0A_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0A_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0A_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0A_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X09_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X09_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0A_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0A_Y0A_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y09_clk_out),
    .clk_out(Tile_X0A_Y0A_clk_out),
    .clk_pass_through(Tile_X0A_Y09_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0A_Y0A_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0A_Y0A_clk_pass_through_out_right),
    .config_config_addr(Tile_X0A_Y09_config_out_config_addr),
    .config_config_data(Tile_X0A_Y09_config_out_config_data),
    .config_out_config_addr(Tile_X0A_Y0A_config_out_config_addr),
    .config_out_config_data(Tile_X0A_Y0A_config_out_config_data),
    .config_out_read(Tile_X0A_Y0A_config_out_read),
    .config_out_write(Tile_X0A_Y0A_config_out_write),
    .config_read(Tile_X0A_Y09_config_out_read),
    .config_write(Tile_X0A_Y09_config_out_write),
    .hi(Tile_X0A_Y0A_hi),
    .lo(Tile_X0A_Y0A_lo_unq1),
    .read_config_data(Tile_X0A_Y0A_read_config_data),
    .read_config_data_in(Tile_X0A_Y09_read_config_data),
    .reset(Tile_X0A_Y09_reset_out),
    .reset_out(Tile_X0A_Y0A_reset_out),
    .stall(Tile_X0A_Y09_stall_out),
    .stall_out(Tile_X0A_Y0A_stall_out),
    .tile_id(Tile_X0A_Y0A_tile_id_in)
);
mantle_wire__typeBit8 Tile_X0A_Y0A_lo (
    .in(Tile_X0A_Y0A_lo_unq1),
    .out(Tile_X0A_Y0A_lo_out)
);
wire [15:0] Tile_X0A_Y0A_tile_id_out;
assign Tile_X0A_Y0A_tile_id_out = {Tile_X0A_Y0A_lo_out[7],Tile_X0A_Y0A_lo_out[7:6],Tile_X0A_Y0A_lo_out[6],Tile_X0A_Y0A_hi[6],Tile_X0A_Y0A_lo_out[5],Tile_X0A_Y0A_hi[5],Tile_X0A_Y0A_lo_out[4:3],Tile_X0A_Y0A_lo_out[3:2],Tile_X0A_Y0A_lo_out[2],Tile_X0A_Y0A_hi[2],Tile_X0A_Y0A_lo_out[1],Tile_X0A_Y0A_hi[1],Tile_X0A_Y0A_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0A_Y0A_tile_id (
    .in(Tile_X0A_Y0A_tile_id_in),
    .out(Tile_X0A_Y0A_tile_id_out)
);
Tile_PE Tile_X0A_Y0B (
    .SB_T0_EAST_SB_IN_B1(Tile_X0B_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0B_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0A_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0A_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0A_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0A_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0A_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0A_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0A_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0A_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0A_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0A_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X09_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X09_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0A_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0A_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0B_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0B_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0A_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0A_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0A_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0A_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0A_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0A_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0A_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0A_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0A_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0A_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X09_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X09_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0A_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0A_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0B_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0B_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0A_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0A_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0A_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0A_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0A_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0A_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0A_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0A_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0A_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0A_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X09_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X09_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0A_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0A_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0B_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0B_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0A_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0A_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0A_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0A_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0A_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0A_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0A_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0A_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0A_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0A_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X09_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X09_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0A_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0A_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0B_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0B_Y0B_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0A_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0A_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0A_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0A_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0A_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0A_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0A_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0A_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0A_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0A_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X09_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X09_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0A_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0A_Y0B_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y0A_clk_out),
    .clk_out(Tile_X0A_Y0B_clk_out),
    .clk_pass_through(Tile_X0A_Y0A_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0A_Y0B_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0A_Y0B_clk_pass_through_out_right),
    .config_config_addr(Tile_X0A_Y0A_config_out_config_addr),
    .config_config_data(Tile_X0A_Y0A_config_out_config_data),
    .config_out_config_addr(Tile_X0A_Y0B_config_out_config_addr),
    .config_out_config_data(Tile_X0A_Y0B_config_out_config_data),
    .config_out_read(Tile_X0A_Y0B_config_out_read),
    .config_out_write(Tile_X0A_Y0B_config_out_write),
    .config_read(Tile_X0A_Y0A_config_out_read),
    .config_write(Tile_X0A_Y0A_config_out_write),
    .hi(Tile_X0A_Y0B_hi_unq1),
    .lo(Tile_X0A_Y0B_lo_unq1),
    .read_config_data(Tile_X0A_Y0B_read_config_data),
    .read_config_data_in(Tile_X0A_Y0A_read_config_data),
    .reset(Tile_X0A_Y0A_reset_out),
    .reset_out(Tile_X0A_Y0B_reset_out),
    .stall(Tile_X0A_Y0A_stall_out),
    .stall_out(Tile_X0A_Y0B_stall_out),
    .tile_id(Tile_X0A_Y0B_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0A_Y0B_hi (
    .in(Tile_X0A_Y0B_hi_unq1),
    .out(Tile_X0A_Y0B_hi_out)
);
mantle_wire__typeBit8 Tile_X0A_Y0B_lo (
    .in(Tile_X0A_Y0B_lo_unq1),
    .out(Tile_X0A_Y0B_lo_out)
);
wire [15:0] Tile_X0A_Y0B_tile_id_out;
assign Tile_X0A_Y0B_tile_id_out = {Tile_X0A_Y0B_lo_out[7],Tile_X0A_Y0B_lo_out[7:6],Tile_X0A_Y0B_lo_out[6],Tile_X0A_Y0B_hi_out[6],Tile_X0A_Y0B_lo_out[5],Tile_X0A_Y0B_hi_out[5],Tile_X0A_Y0B_lo_out[4:3],Tile_X0A_Y0B_lo_out[3:2],Tile_X0A_Y0B_lo_out[2],Tile_X0A_Y0B_hi_out[2],Tile_X0A_Y0B_lo_out[1],Tile_X0A_Y0B_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X0A_Y0B_tile_id (
    .in(Tile_X0A_Y0B_tile_id_in),
    .out(Tile_X0A_Y0B_tile_id_out)
);
Tile_PE Tile_X0A_Y0C (
    .SB_T0_EAST_SB_IN_B1(Tile_X0B_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0B_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0A_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0A_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0A_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0A_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0A_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0A_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0A_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0A_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0A_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0A_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X09_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X09_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0A_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0A_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0B_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0B_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0A_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0A_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0A_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0A_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0A_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0A_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0A_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0A_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0A_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0A_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X09_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X09_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0A_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0A_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0B_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0B_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0A_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0A_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0A_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0A_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0A_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0A_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0A_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0A_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0A_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0A_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X09_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X09_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0A_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0A_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0B_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0B_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0A_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0A_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0A_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0A_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0A_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0A_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0A_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0A_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0A_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0A_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X09_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X09_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0A_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0A_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0B_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0B_Y0C_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0A_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0A_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0A_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0A_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0A_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0A_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0A_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0A_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0A_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0A_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X09_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X09_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0A_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0A_Y0C_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y0B_clk_out),
    .clk_out(Tile_X0A_Y0C_clk_out),
    .clk_pass_through(Tile_X0A_Y0B_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0A_Y0C_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0A_Y0C_clk_pass_through_out_right),
    .config_config_addr(Tile_X0A_Y0B_config_out_config_addr),
    .config_config_data(Tile_X0A_Y0B_config_out_config_data),
    .config_out_config_addr(Tile_X0A_Y0C_config_out_config_addr),
    .config_out_config_data(Tile_X0A_Y0C_config_out_config_data),
    .config_out_read(Tile_X0A_Y0C_config_out_read),
    .config_out_write(Tile_X0A_Y0C_config_out_write),
    .config_read(Tile_X0A_Y0B_config_out_read),
    .config_write(Tile_X0A_Y0B_config_out_write),
    .hi(Tile_X0A_Y0C_hi_unq1),
    .lo(Tile_X0A_Y0C_lo_unq1),
    .read_config_data(Tile_X0A_Y0C_read_config_data),
    .read_config_data_in(Tile_X0A_Y0B_read_config_data),
    .reset(Tile_X0A_Y0B_reset_out),
    .reset_out(Tile_X0A_Y0C_reset_out),
    .stall(Tile_X0A_Y0B_stall_out),
    .stall_out(Tile_X0A_Y0C_stall_out),
    .tile_id(Tile_X0A_Y0C_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0A_Y0C_hi (
    .in(Tile_X0A_Y0C_hi_unq1),
    .out(Tile_X0A_Y0C_hi_out)
);
mantle_wire__typeBit8 Tile_X0A_Y0C_lo (
    .in(Tile_X0A_Y0C_lo_unq1),
    .out(Tile_X0A_Y0C_lo_out)
);
wire [15:0] Tile_X0A_Y0C_tile_id_out;
assign Tile_X0A_Y0C_tile_id_out = {Tile_X0A_Y0C_lo_out[7],Tile_X0A_Y0C_lo_out[7:6],Tile_X0A_Y0C_lo_out[6],Tile_X0A_Y0C_hi_out[6],Tile_X0A_Y0C_lo_out[5],Tile_X0A_Y0C_hi_out[5],Tile_X0A_Y0C_lo_out[4:3],Tile_X0A_Y0C_lo_out[3:2],Tile_X0A_Y0C_lo_out[2],Tile_X0A_Y0C_hi_out[2:1],Tile_X0A_Y0C_lo_out[0],Tile_X0A_Y0C_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0A_Y0C_tile_id (
    .in(Tile_X0A_Y0C_tile_id_in),
    .out(Tile_X0A_Y0C_tile_id_out)
);
Tile_PE Tile_X0A_Y0D (
    .SB_T0_EAST_SB_IN_B1(Tile_X0B_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0B_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0A_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0A_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0A_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0A_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0A_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0A_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0A_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0A_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0A_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0A_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X09_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X09_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0A_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0A_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0B_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0B_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0A_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0A_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0A_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0A_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0A_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0A_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0A_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0A_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0A_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0A_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X09_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X09_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0A_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0A_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0B_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0B_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0A_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0A_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0A_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0A_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0A_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0A_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0A_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0A_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0A_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0A_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X09_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X09_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0A_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0A_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0B_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0B_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0A_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0A_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0A_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0A_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0A_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0A_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0A_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0A_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0A_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0A_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X09_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X09_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0A_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0A_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0B_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0B_Y0D_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0A_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0A_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0A_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0A_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0A_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0A_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0A_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0A_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0A_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0A_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X09_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X09_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0A_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0A_Y0D_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y0C_clk_out),
    .clk_out(Tile_X0A_Y0D_clk_out),
    .clk_pass_through(Tile_X0A_Y0C_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0A_Y0D_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0A_Y0D_clk_pass_through_out_right),
    .config_config_addr(Tile_X0A_Y0C_config_out_config_addr),
    .config_config_data(Tile_X0A_Y0C_config_out_config_data),
    .config_out_config_addr(Tile_X0A_Y0D_config_out_config_addr),
    .config_out_config_data(Tile_X0A_Y0D_config_out_config_data),
    .config_out_read(Tile_X0A_Y0D_config_out_read),
    .config_out_write(Tile_X0A_Y0D_config_out_write),
    .config_read(Tile_X0A_Y0C_config_out_read),
    .config_write(Tile_X0A_Y0C_config_out_write),
    .hi(Tile_X0A_Y0D_hi_unq1),
    .lo(Tile_X0A_Y0D_lo_unq1),
    .read_config_data(Tile_X0A_Y0D_read_config_data),
    .read_config_data_in(Tile_X0A_Y0C_read_config_data),
    .reset(Tile_X0A_Y0C_reset_out),
    .reset_out(Tile_X0A_Y0D_reset_out),
    .stall(Tile_X0A_Y0C_stall_out),
    .stall_out(Tile_X0A_Y0D_stall_out),
    .tile_id(Tile_X0A_Y0D_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0A_Y0D_hi (
    .in(Tile_X0A_Y0D_hi_unq1),
    .out(Tile_X0A_Y0D_hi_out)
);
mantle_wire__typeBit8 Tile_X0A_Y0D_lo (
    .in(Tile_X0A_Y0D_lo_unq1),
    .out(Tile_X0A_Y0D_lo_out)
);
wire [15:0] Tile_X0A_Y0D_tile_id_out;
assign Tile_X0A_Y0D_tile_id_out = {Tile_X0A_Y0D_lo_out[7],Tile_X0A_Y0D_lo_out[7:6],Tile_X0A_Y0D_lo_out[6],Tile_X0A_Y0D_hi_out[6],Tile_X0A_Y0D_lo_out[5],Tile_X0A_Y0D_hi_out[5],Tile_X0A_Y0D_lo_out[4:3],Tile_X0A_Y0D_lo_out[3:2],Tile_X0A_Y0D_lo_out[2],Tile_X0A_Y0D_hi_out[2:1],Tile_X0A_Y0D_lo_out[0],Tile_X0A_Y0D_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X0A_Y0D_tile_id (
    .in(Tile_X0A_Y0D_tile_id_in),
    .out(Tile_X0A_Y0D_tile_id_out)
);
Tile_PE Tile_X0A_Y0E (
    .SB_T0_EAST_SB_IN_B1(Tile_X0B_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0B_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0A_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0A_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0A_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0A_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0A_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0A_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0A_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0A_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0A_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0A_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X09_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X09_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0A_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0A_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0B_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0B_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0A_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0A_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0A_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0A_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0A_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0A_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0A_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0A_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0A_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0A_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X09_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X09_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0A_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0A_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0B_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0B_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0A_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0A_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0A_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0A_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0A_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0A_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0A_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0A_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0A_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0A_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X09_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X09_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0A_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0A_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0B_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0B_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0A_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0A_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0A_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0A_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0A_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0A_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0A_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0A_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0A_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0A_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X09_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X09_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0A_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0A_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0B_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0B_Y0E_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0A_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0A_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0A_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0A_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0A_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0A_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0A_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0A_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0A_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0A_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X09_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X09_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0A_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0A_Y0E_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y0D_clk_out),
    .clk_out(Tile_X0A_Y0E_clk_out),
    .clk_pass_through(Tile_X0A_Y0D_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0A_Y0E_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0A_Y0E_clk_pass_through_out_right),
    .config_config_addr(Tile_X0A_Y0D_config_out_config_addr),
    .config_config_data(Tile_X0A_Y0D_config_out_config_data),
    .config_out_config_addr(Tile_X0A_Y0E_config_out_config_addr),
    .config_out_config_data(Tile_X0A_Y0E_config_out_config_data),
    .config_out_read(Tile_X0A_Y0E_config_out_read),
    .config_out_write(Tile_X0A_Y0E_config_out_write),
    .config_read(Tile_X0A_Y0D_config_out_read),
    .config_write(Tile_X0A_Y0D_config_out_write),
    .hi(Tile_X0A_Y0E_hi_unq1),
    .lo(Tile_X0A_Y0E_lo_unq1),
    .read_config_data(Tile_X0A_Y0E_read_config_data),
    .read_config_data_in(Tile_X0A_Y0D_read_config_data),
    .reset(Tile_X0A_Y0D_reset_out),
    .reset_out(Tile_X0A_Y0E_reset_out),
    .stall(Tile_X0A_Y0D_stall_out),
    .stall_out(Tile_X0A_Y0E_stall_out),
    .tile_id(Tile_X0A_Y0E_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0A_Y0E_hi (
    .in(Tile_X0A_Y0E_hi_unq1),
    .out(Tile_X0A_Y0E_hi_out)
);
mantle_wire__typeBit8 Tile_X0A_Y0E_lo (
    .in(Tile_X0A_Y0E_lo_unq1),
    .out(Tile_X0A_Y0E_lo_out)
);
wire [15:0] Tile_X0A_Y0E_tile_id_out;
assign Tile_X0A_Y0E_tile_id_out = {Tile_X0A_Y0E_lo_out[7],Tile_X0A_Y0E_lo_out[7:6],Tile_X0A_Y0E_lo_out[6],Tile_X0A_Y0E_hi_out[6],Tile_X0A_Y0E_lo_out[5],Tile_X0A_Y0E_hi_out[5],Tile_X0A_Y0E_lo_out[4:3],Tile_X0A_Y0E_lo_out[3:2],Tile_X0A_Y0E_lo_out[2],Tile_X0A_Y0E_hi_out[2:1],Tile_X0A_Y0E_hi_out[1],Tile_X0A_Y0E_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0A_Y0E_tile_id (
    .in(Tile_X0A_Y0E_tile_id_in),
    .out(Tile_X0A_Y0E_tile_id_out)
);
Tile_PE Tile_X0A_Y0F (
    .SB_T0_EAST_SB_IN_B1(Tile_X0B_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0B_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0A_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0A_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0A_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0A_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0A_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0A_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0A_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0A_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0A_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0A_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X09_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X09_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0A_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0A_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0B_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0B_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0A_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0A_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0A_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0A_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0A_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0A_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0A_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0A_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0A_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0A_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X09_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X09_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0A_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0A_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0B_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0B_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0A_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0A_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0A_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0A_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0A_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0A_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0A_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0A_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0A_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0A_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X09_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X09_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0A_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0A_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0B_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0B_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0A_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0A_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0A_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0A_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0A_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0A_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0A_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0A_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0A_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0A_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X09_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X09_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0A_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0A_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0B_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0B_Y0F_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0A_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0A_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0A_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0A_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0A_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0A_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0A_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0A_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0A_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0A_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X09_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X09_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0A_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0A_Y0F_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y0E_clk_out),
    .clk_out(Tile_X0A_Y0F_clk_out),
    .clk_pass_through(Tile_X0A_Y0E_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0A_Y0F_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0A_Y0F_clk_pass_through_out_right),
    .config_config_addr(Tile_X0A_Y0E_config_out_config_addr),
    .config_config_data(Tile_X0A_Y0E_config_out_config_data),
    .config_out_config_addr(Tile_X0A_Y0F_config_out_config_addr),
    .config_out_config_data(Tile_X0A_Y0F_config_out_config_data),
    .config_out_read(Tile_X0A_Y0F_config_out_read),
    .config_out_write(Tile_X0A_Y0F_config_out_write),
    .config_read(Tile_X0A_Y0E_config_out_read),
    .config_write(Tile_X0A_Y0E_config_out_write),
    .hi(Tile_X0A_Y0F_hi_unq1),
    .lo(Tile_X0A_Y0F_lo_unq1),
    .read_config_data(Tile_X0A_Y0F_read_config_data),
    .read_config_data_in(Tile_X0A_Y0E_read_config_data),
    .reset(Tile_X0A_Y0E_reset_out),
    .reset_out(Tile_X0A_Y0F_reset_out),
    .stall(Tile_X0A_Y0E_stall_out),
    .stall_out(Tile_X0A_Y0F_stall_out),
    .tile_id(Tile_X0A_Y0F_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0A_Y0F_hi (
    .in(Tile_X0A_Y0F_hi_unq1),
    .out(Tile_X0A_Y0F_hi_out)
);
mantle_wire__typeBit8 Tile_X0A_Y0F_lo (
    .in(Tile_X0A_Y0F_lo_unq1),
    .out(Tile_X0A_Y0F_lo_out)
);
wire [15:0] Tile_X0A_Y0F_tile_id_out;
assign Tile_X0A_Y0F_tile_id_out = {Tile_X0A_Y0F_lo_out[7],Tile_X0A_Y0F_lo_out[7:6],Tile_X0A_Y0F_lo_out[6],Tile_X0A_Y0F_hi_out[6],Tile_X0A_Y0F_lo_out[5],Tile_X0A_Y0F_hi_out[5],Tile_X0A_Y0F_lo_out[4:3],Tile_X0A_Y0F_lo_out[3:2],Tile_X0A_Y0F_lo_out[2],Tile_X0A_Y0F_hi_out[2:1],Tile_X0A_Y0F_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X0A_Y0F_tile_id (
    .in(Tile_X0A_Y0F_tile_id_in),
    .out(Tile_X0A_Y0F_tile_id_out)
);
Tile_PE Tile_X0A_Y10 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0B_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0B_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0A_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0A_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0A_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0A_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0A_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0A_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T0_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0A_Y10_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0A_Y10_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X09_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X09_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0A_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0A_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0B_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0B_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0A_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0A_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0A_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0A_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0A_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0A_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T1_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0A_Y10_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0A_Y10_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X09_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X09_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0A_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0A_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0B_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0B_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0A_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0A_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0A_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0A_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0A_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0A_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T2_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0A_Y10_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0A_Y10_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X09_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X09_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0A_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0A_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0B_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0B_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0A_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0A_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0A_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0A_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0A_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0A_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T3_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0A_Y10_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0A_Y10_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X09_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X09_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0A_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0A_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0B_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0B_Y10_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0A_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0A_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0A_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0A_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0A_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0A_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T4_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0A_Y10_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0A_Y10_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X09_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X09_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0A_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0A_Y10_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y0F_clk_out),
    .clk_out(Tile_X0A_Y10_clk_out),
    .clk_pass_through(Tile_X0A_Y0F_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0A_Y10_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0A_Y10_clk_pass_through_out_right),
    .config_config_addr(Tile_X0A_Y0F_config_out_config_addr),
    .config_config_data(Tile_X0A_Y0F_config_out_config_data),
    .config_out_config_addr(Tile_X0A_Y10_config_out_config_addr),
    .config_out_config_data(Tile_X0A_Y10_config_out_config_data),
    .config_out_read(Tile_X0A_Y10_config_out_read),
    .config_out_write(Tile_X0A_Y10_config_out_write),
    .config_read(Tile_X0A_Y0F_config_out_read),
    .config_write(Tile_X0A_Y0F_config_out_write),
    .hi(Tile_X0A_Y10_hi),
    .lo(Tile_X0A_Y10_lo_unq1),
    .read_config_data(Tile_X0A_Y10_read_config_data),
    .read_config_data_in(Tile_X0A_Y0F_read_config_data),
    .reset(Tile_X0A_Y0F_reset_out),
    .reset_out(Tile_X0A_Y10_reset_out),
    .stall(Tile_X0A_Y0F_stall_out),
    .stall_out(Tile_X0A_Y10_stall_out),
    .tile_id(Tile_X0A_Y10_tile_id_in)
);
mantle_wire__typeBit8 Tile_X0A_Y10_lo (
    .in(Tile_X0A_Y10_lo_unq1),
    .out(Tile_X0A_Y10_lo_out)
);
wire [15:0] Tile_X0A_Y10_tile_id_out;
assign Tile_X0A_Y10_tile_id_out = {Tile_X0A_Y10_lo_out[7],Tile_X0A_Y10_lo_out[7:6],Tile_X0A_Y10_lo_out[6],Tile_X0A_Y10_hi[6],Tile_X0A_Y10_lo_out[5],Tile_X0A_Y10_hi[5],Tile_X0A_Y10_lo_out[4:3],Tile_X0A_Y10_lo_out[3:2],Tile_X0A_Y10_hi[2],Tile_X0A_Y10_lo_out[1],Tile_X0A_Y10_lo_out[1:0],Tile_X0A_Y10_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0A_Y10_tile_id (
    .in(Tile_X0A_Y10_tile_id_in),
    .out(Tile_X0A_Y10_tile_id_out)
);
wire [15:0] Tile_X0B_Y00_tile_id;
assign Tile_X0B_Y00_tile_id = {Tile_X0B_Y00_lo[7],Tile_X0B_Y00_lo[7:6],Tile_X0B_Y00_lo[6],Tile_X0B_Y00_hi[6],Tile_X0B_Y00_lo[5],Tile_X0B_Y00_hi[5:4],Tile_X0B_Y00_lo[3],Tile_X0B_Y00_lo[3:2],Tile_X0B_Y00_lo[2:1],Tile_X0B_Y00_lo[1:0],Tile_X0B_Y00_lo[0]};
Tile_io_core Tile_X0B_Y00 (
    .tile_id(Tile_X0B_Y00_tile_id),
    .glb2io_1(glb2io_1_X0B_Y00),
    .f2io_1(Tile_X0B_Y01_SB_T0_NORTH_SB_OUT_B1),
    .io2glb_1(Tile_X0B_Y00_io2glb_1),
    .io2f_1(Tile_X0B_Y00_io2f_1),
    .glb2io_16(glb2io_16_X0B_Y00),
    .f2io_16(Tile_X0B_Y01_SB_T0_NORTH_SB_OUT_B16),
    .io2glb_16(Tile_X0B_Y00_io2glb_16),
    .io2f_16(Tile_X0B_Y00_io2f_16),
    .hi(Tile_X0B_Y00_hi),
    .lo(Tile_X0B_Y00_lo)
);
Tile_MemCore Tile_X0B_Y01 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0C_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0C_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0B_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0B_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0B_Y00_io2f_1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0B_Y00_io2f_16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0B_Y01_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0B_Y01_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0B_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0B_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0B_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0B_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0A_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0A_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0B_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0B_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0C_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0C_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0B_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0B_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0B_Y00_io2f_1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0B_Y00_io2f_16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0B_Y01_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0B_Y01_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0B_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0B_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0B_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0B_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0A_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0A_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0B_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0B_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0C_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0C_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0B_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0B_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0B_Y00_io2f_1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0B_Y00_io2f_16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0B_Y01_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0B_Y01_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0B_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0B_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0B_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0B_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0A_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0A_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0B_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0B_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0C_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0C_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0B_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0B_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0B_Y00_io2f_1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0B_Y00_io2f_16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0B_Y01_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0B_Y01_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0B_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0B_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0B_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0B_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0A_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0A_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0B_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0B_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0C_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0C_Y01_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0B_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0B_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0B_Y00_io2f_1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0B_Y00_io2f_16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0B_Y01_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0B_Y01_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0B_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0B_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0B_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0B_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0A_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0A_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0B_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0B_Y01_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y01_clk_pass_through_out_right),
    .clk_out(Tile_X0B_Y01_clk_out),
    .config_config_addr(config_11_config_addr),
    .config_config_data(config_11_config_data),
    .config_out_config_addr(Tile_X0B_Y01_config_out_config_addr),
    .config_out_config_data(Tile_X0B_Y01_config_out_config_data),
    .config_out_read(Tile_X0B_Y01_config_out_read),
    .config_out_write(Tile_X0B_Y01_config_out_write),
    .config_read(config_11_read),
    .config_write(config_11_write),
    .hi(Tile_X0B_Y01_hi_unq1),
    .lo(Tile_X0B_Y01_lo_unq1),
    .read_config_data(Tile_X0B_Y01_read_config_data),
    .read_config_data_in(const_0_32_out),
    .reset(reset),
    .reset_out(Tile_X0B_Y01_reset_out),
    .stall(stall[11]),
    .stall_out(Tile_X0B_Y01_stall_out),
    .tile_id(Tile_X0B_Y01_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0B_Y01_hi (
    .in(Tile_X0B_Y01_hi_unq1),
    .out(Tile_X0B_Y01_hi_out)
);
mantle_wire__typeBit8 Tile_X0B_Y01_lo (
    .in(Tile_X0B_Y01_lo_unq1),
    .out(Tile_X0B_Y01_lo_out)
);
wire [15:0] Tile_X0B_Y01_tile_id_out;
assign Tile_X0B_Y01_tile_id_out = {Tile_X0B_Y01_lo_out[7],Tile_X0B_Y01_lo_out[7:6],Tile_X0B_Y01_lo_out[6],Tile_X0B_Y01_hi_out[6],Tile_X0B_Y01_lo_out[5],Tile_X0B_Y01_hi_out[5:4],Tile_X0B_Y01_lo_out[3],Tile_X0B_Y01_lo_out[3:2],Tile_X0B_Y01_lo_out[2:1],Tile_X0B_Y01_lo_out[1:0],Tile_X0B_Y01_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X0B_Y01_tile_id (
    .in(Tile_X0B_Y01_tile_id_in),
    .out(Tile_X0B_Y01_tile_id_out)
);
Tile_MemCore Tile_X0B_Y02 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0C_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0C_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0B_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0B_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0B_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0B_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0B_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0B_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0B_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0B_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0B_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0B_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0A_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0A_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0B_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0B_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0C_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0C_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0B_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0B_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0B_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0B_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0B_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0B_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0B_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0B_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0B_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0B_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0A_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0A_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0B_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0B_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0C_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0C_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0B_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0B_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0B_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0B_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0B_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0B_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0B_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0B_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0B_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0B_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0A_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0A_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0B_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0B_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0C_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0C_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0B_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0B_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0B_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0B_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0B_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0B_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0B_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0B_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0B_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0B_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0A_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0A_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0B_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0B_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0C_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0C_Y02_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0B_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0B_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0B_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0B_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0B_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0B_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0B_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0B_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0B_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0B_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0A_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0A_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0B_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0B_Y02_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y02_clk_pass_through_out_right),
    .clk_out(Tile_X0B_Y02_clk_out),
    .config_config_addr(Tile_X0B_Y01_config_out_config_addr),
    .config_config_data(Tile_X0B_Y01_config_out_config_data),
    .config_out_config_addr(Tile_X0B_Y02_config_out_config_addr),
    .config_out_config_data(Tile_X0B_Y02_config_out_config_data),
    .config_out_read(Tile_X0B_Y02_config_out_read),
    .config_out_write(Tile_X0B_Y02_config_out_write),
    .config_read(Tile_X0B_Y01_config_out_read),
    .config_write(Tile_X0B_Y01_config_out_write),
    .hi(Tile_X0B_Y02_hi_unq1),
    .lo(Tile_X0B_Y02_lo_unq1),
    .read_config_data(Tile_X0B_Y02_read_config_data),
    .read_config_data_in(Tile_X0B_Y01_read_config_data),
    .reset(Tile_X0B_Y01_reset_out),
    .reset_out(Tile_X0B_Y02_reset_out),
    .stall(Tile_X0B_Y01_stall_out),
    .stall_out(Tile_X0B_Y02_stall_out),
    .tile_id(Tile_X0B_Y02_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0B_Y02_hi (
    .in(Tile_X0B_Y02_hi_unq1),
    .out(Tile_X0B_Y02_hi_out)
);
mantle_wire__typeBit8 Tile_X0B_Y02_lo (
    .in(Tile_X0B_Y02_lo_unq1),
    .out(Tile_X0B_Y02_lo_out)
);
wire [15:0] Tile_X0B_Y02_tile_id_out;
assign Tile_X0B_Y02_tile_id_out = {Tile_X0B_Y02_lo_out[7],Tile_X0B_Y02_lo_out[7:6],Tile_X0B_Y02_lo_out[6],Tile_X0B_Y02_hi_out[6],Tile_X0B_Y02_lo_out[5],Tile_X0B_Y02_hi_out[5:4],Tile_X0B_Y02_lo_out[3],Tile_X0B_Y02_lo_out[3:2],Tile_X0B_Y02_lo_out[2:1],Tile_X0B_Y02_lo_out[1],Tile_X0B_Y02_hi_out[1],Tile_X0B_Y02_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0B_Y02_tile_id (
    .in(Tile_X0B_Y02_tile_id_in),
    .out(Tile_X0B_Y02_tile_id_out)
);
Tile_MemCore Tile_X0B_Y03 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0C_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0C_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0B_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0B_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0B_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0B_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0B_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0B_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0B_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0B_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0B_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0B_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0A_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0A_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0B_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0B_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0C_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0C_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0B_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0B_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0B_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0B_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0B_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0B_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0B_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0B_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0B_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0B_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0A_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0A_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0B_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0B_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0C_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0C_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0B_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0B_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0B_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0B_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0B_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0B_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0B_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0B_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0B_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0B_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0A_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0A_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0B_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0B_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0C_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0C_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0B_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0B_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0B_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0B_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0B_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0B_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0B_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0B_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0B_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0B_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0A_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0A_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0B_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0B_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0C_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0C_Y03_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0B_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0B_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0B_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0B_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0B_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0B_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0B_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0B_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0B_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0B_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0A_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0A_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0B_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0B_Y03_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y03_clk_pass_through_out_right),
    .clk_out(Tile_X0B_Y03_clk_out),
    .config_config_addr(Tile_X0B_Y02_config_out_config_addr),
    .config_config_data(Tile_X0B_Y02_config_out_config_data),
    .config_out_config_addr(Tile_X0B_Y03_config_out_config_addr),
    .config_out_config_data(Tile_X0B_Y03_config_out_config_data),
    .config_out_read(Tile_X0B_Y03_config_out_read),
    .config_out_write(Tile_X0B_Y03_config_out_write),
    .config_read(Tile_X0B_Y02_config_out_read),
    .config_write(Tile_X0B_Y02_config_out_write),
    .hi(Tile_X0B_Y03_hi_unq1),
    .lo(Tile_X0B_Y03_lo_unq1),
    .read_config_data(Tile_X0B_Y03_read_config_data),
    .read_config_data_in(Tile_X0B_Y02_read_config_data),
    .reset(Tile_X0B_Y02_reset_out),
    .reset_out(Tile_X0B_Y03_reset_out),
    .stall(Tile_X0B_Y02_stall_out),
    .stall_out(Tile_X0B_Y03_stall_out),
    .tile_id(Tile_X0B_Y03_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0B_Y03_hi (
    .in(Tile_X0B_Y03_hi_unq1),
    .out(Tile_X0B_Y03_hi_out)
);
mantle_wire__typeBit8 Tile_X0B_Y03_lo (
    .in(Tile_X0B_Y03_lo_unq1),
    .out(Tile_X0B_Y03_lo_out)
);
wire [15:0] Tile_X0B_Y03_tile_id_out;
assign Tile_X0B_Y03_tile_id_out = {Tile_X0B_Y03_lo_out[7],Tile_X0B_Y03_lo_out[7:6],Tile_X0B_Y03_lo_out[6],Tile_X0B_Y03_hi_out[6],Tile_X0B_Y03_lo_out[5],Tile_X0B_Y03_hi_out[5:4],Tile_X0B_Y03_lo_out[3],Tile_X0B_Y03_lo_out[3:2],Tile_X0B_Y03_lo_out[2:1],Tile_X0B_Y03_lo_out[1],Tile_X0B_Y03_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X0B_Y03_tile_id (
    .in(Tile_X0B_Y03_tile_id_in),
    .out(Tile_X0B_Y03_tile_id_out)
);
Tile_MemCore Tile_X0B_Y04 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0C_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0C_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0B_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0B_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0B_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0B_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0B_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0B_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0B_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0B_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0B_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0B_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0A_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0A_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0B_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0B_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0C_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0C_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0B_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0B_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0B_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0B_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0B_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0B_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0B_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0B_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0B_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0B_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0A_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0A_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0B_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0B_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0C_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0C_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0B_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0B_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0B_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0B_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0B_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0B_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0B_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0B_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0B_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0B_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0A_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0A_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0B_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0B_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0C_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0C_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0B_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0B_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0B_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0B_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0B_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0B_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0B_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0B_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0B_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0B_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0A_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0A_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0B_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0B_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0C_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0C_Y04_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0B_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0B_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0B_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0B_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0B_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0B_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0B_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0B_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0B_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0B_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0A_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0A_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0B_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0B_Y04_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y04_clk_pass_through_out_right),
    .clk_out(Tile_X0B_Y04_clk_out),
    .config_config_addr(Tile_X0B_Y03_config_out_config_addr),
    .config_config_data(Tile_X0B_Y03_config_out_config_data),
    .config_out_config_addr(Tile_X0B_Y04_config_out_config_addr),
    .config_out_config_data(Tile_X0B_Y04_config_out_config_data),
    .config_out_read(Tile_X0B_Y04_config_out_read),
    .config_out_write(Tile_X0B_Y04_config_out_write),
    .config_read(Tile_X0B_Y03_config_out_read),
    .config_write(Tile_X0B_Y03_config_out_write),
    .hi(Tile_X0B_Y04_hi_unq1),
    .lo(Tile_X0B_Y04_lo_unq1),
    .read_config_data(Tile_X0B_Y04_read_config_data),
    .read_config_data_in(Tile_X0B_Y03_read_config_data),
    .reset(Tile_X0B_Y03_reset_out),
    .reset_out(Tile_X0B_Y04_reset_out),
    .stall(Tile_X0B_Y03_stall_out),
    .stall_out(Tile_X0B_Y04_stall_out),
    .tile_id(Tile_X0B_Y04_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0B_Y04_hi (
    .in(Tile_X0B_Y04_hi_unq1),
    .out(Tile_X0B_Y04_hi_out)
);
mantle_wire__typeBit8 Tile_X0B_Y04_lo (
    .in(Tile_X0B_Y04_lo_unq1),
    .out(Tile_X0B_Y04_lo_out)
);
wire [15:0] Tile_X0B_Y04_tile_id_out;
assign Tile_X0B_Y04_tile_id_out = {Tile_X0B_Y04_lo_out[7],Tile_X0B_Y04_lo_out[7:6],Tile_X0B_Y04_lo_out[6],Tile_X0B_Y04_hi_out[6],Tile_X0B_Y04_lo_out[5],Tile_X0B_Y04_hi_out[5:4],Tile_X0B_Y04_lo_out[3],Tile_X0B_Y04_lo_out[3:2],Tile_X0B_Y04_lo_out[2:1],Tile_X0B_Y04_hi_out[1],Tile_X0B_Y04_lo_out[0],Tile_X0B_Y04_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0B_Y04_tile_id (
    .in(Tile_X0B_Y04_tile_id_in),
    .out(Tile_X0B_Y04_tile_id_out)
);
Tile_MemCore Tile_X0B_Y05 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0C_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0C_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0B_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0B_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0B_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0B_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0B_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0B_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0B_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0B_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0B_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0B_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0A_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0A_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0B_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0B_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0C_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0C_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0B_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0B_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0B_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0B_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0B_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0B_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0B_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0B_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0B_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0B_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0A_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0A_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0B_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0B_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0C_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0C_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0B_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0B_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0B_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0B_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0B_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0B_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0B_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0B_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0B_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0B_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0A_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0A_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0B_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0B_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0C_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0C_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0B_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0B_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0B_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0B_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0B_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0B_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0B_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0B_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0B_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0B_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0A_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0A_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0B_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0B_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0C_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0C_Y05_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0B_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0B_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0B_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0B_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0B_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0B_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0B_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0B_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0B_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0B_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0A_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0A_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0B_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0B_Y05_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y05_clk_pass_through_out_right),
    .clk_out(Tile_X0B_Y05_clk_out),
    .config_config_addr(Tile_X0B_Y04_config_out_config_addr),
    .config_config_data(Tile_X0B_Y04_config_out_config_data),
    .config_out_config_addr(Tile_X0B_Y05_config_out_config_addr),
    .config_out_config_data(Tile_X0B_Y05_config_out_config_data),
    .config_out_read(Tile_X0B_Y05_config_out_read),
    .config_out_write(Tile_X0B_Y05_config_out_write),
    .config_read(Tile_X0B_Y04_config_out_read),
    .config_write(Tile_X0B_Y04_config_out_write),
    .hi(Tile_X0B_Y05_hi_unq1),
    .lo(Tile_X0B_Y05_lo_unq1),
    .read_config_data(Tile_X0B_Y05_read_config_data),
    .read_config_data_in(Tile_X0B_Y04_read_config_data),
    .reset(Tile_X0B_Y04_reset_out),
    .reset_out(Tile_X0B_Y05_reset_out),
    .stall(Tile_X0B_Y04_stall_out),
    .stall_out(Tile_X0B_Y05_stall_out),
    .tile_id(Tile_X0B_Y05_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0B_Y05_hi (
    .in(Tile_X0B_Y05_hi_unq1),
    .out(Tile_X0B_Y05_hi_out)
);
mantle_wire__typeBit8 Tile_X0B_Y05_lo (
    .in(Tile_X0B_Y05_lo_unq1),
    .out(Tile_X0B_Y05_lo_out)
);
wire [15:0] Tile_X0B_Y05_tile_id_out;
assign Tile_X0B_Y05_tile_id_out = {Tile_X0B_Y05_lo_out[7],Tile_X0B_Y05_lo_out[7:6],Tile_X0B_Y05_lo_out[6],Tile_X0B_Y05_hi_out[6],Tile_X0B_Y05_lo_out[5],Tile_X0B_Y05_hi_out[5:4],Tile_X0B_Y05_lo_out[3],Tile_X0B_Y05_lo_out[3:2],Tile_X0B_Y05_lo_out[2:1],Tile_X0B_Y05_hi_out[1],Tile_X0B_Y05_lo_out[0],Tile_X0B_Y05_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X0B_Y05_tile_id (
    .in(Tile_X0B_Y05_tile_id_in),
    .out(Tile_X0B_Y05_tile_id_out)
);
Tile_MemCore Tile_X0B_Y06 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0C_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0C_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0B_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0B_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0B_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0B_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0B_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0B_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0B_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0B_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0B_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0B_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0A_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0A_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0B_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0B_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0C_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0C_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0B_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0B_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0B_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0B_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0B_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0B_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0B_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0B_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0B_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0B_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0A_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0A_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0B_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0B_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0C_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0C_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0B_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0B_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0B_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0B_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0B_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0B_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0B_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0B_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0B_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0B_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0A_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0A_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0B_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0B_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0C_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0C_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0B_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0B_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0B_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0B_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0B_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0B_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0B_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0B_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0B_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0B_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0A_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0A_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0B_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0B_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0C_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0C_Y06_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0B_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0B_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0B_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0B_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0B_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0B_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0B_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0B_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0B_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0B_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0A_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0A_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0B_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0B_Y06_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y06_clk_pass_through_out_right),
    .clk_out(Tile_X0B_Y06_clk_out),
    .config_config_addr(Tile_X0B_Y05_config_out_config_addr),
    .config_config_data(Tile_X0B_Y05_config_out_config_data),
    .config_out_config_addr(Tile_X0B_Y06_config_out_config_addr),
    .config_out_config_data(Tile_X0B_Y06_config_out_config_data),
    .config_out_read(Tile_X0B_Y06_config_out_read),
    .config_out_write(Tile_X0B_Y06_config_out_write),
    .config_read(Tile_X0B_Y05_config_out_read),
    .config_write(Tile_X0B_Y05_config_out_write),
    .hi(Tile_X0B_Y06_hi_unq1),
    .lo(Tile_X0B_Y06_lo_unq1),
    .read_config_data(Tile_X0B_Y06_read_config_data),
    .read_config_data_in(Tile_X0B_Y05_read_config_data),
    .reset(Tile_X0B_Y05_reset_out),
    .reset_out(Tile_X0B_Y06_reset_out),
    .stall(Tile_X0B_Y05_stall_out),
    .stall_out(Tile_X0B_Y06_stall_out),
    .tile_id(Tile_X0B_Y06_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0B_Y06_hi (
    .in(Tile_X0B_Y06_hi_unq1),
    .out(Tile_X0B_Y06_hi_out)
);
mantle_wire__typeBit8 Tile_X0B_Y06_lo (
    .in(Tile_X0B_Y06_lo_unq1),
    .out(Tile_X0B_Y06_lo_out)
);
wire [15:0] Tile_X0B_Y06_tile_id_out;
assign Tile_X0B_Y06_tile_id_out = {Tile_X0B_Y06_lo_out[7],Tile_X0B_Y06_lo_out[7:6],Tile_X0B_Y06_lo_out[6],Tile_X0B_Y06_hi_out[6],Tile_X0B_Y06_lo_out[5],Tile_X0B_Y06_hi_out[5:4],Tile_X0B_Y06_lo_out[3],Tile_X0B_Y06_lo_out[3:2],Tile_X0B_Y06_lo_out[2:1],Tile_X0B_Y06_hi_out[1],Tile_X0B_Y06_hi_out[1],Tile_X0B_Y06_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0B_Y06_tile_id (
    .in(Tile_X0B_Y06_tile_id_in),
    .out(Tile_X0B_Y06_tile_id_out)
);
Tile_MemCore Tile_X0B_Y07 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0C_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0C_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0B_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0B_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0B_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0B_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0B_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0B_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0B_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0B_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0B_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0B_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0A_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0A_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0B_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0B_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0C_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0C_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0B_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0B_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0B_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0B_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0B_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0B_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0B_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0B_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0B_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0B_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0A_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0A_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0B_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0B_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0C_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0C_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0B_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0B_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0B_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0B_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0B_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0B_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0B_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0B_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0B_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0B_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0A_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0A_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0B_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0B_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0C_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0C_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0B_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0B_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0B_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0B_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0B_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0B_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0B_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0B_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0B_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0B_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0A_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0A_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0B_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0B_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0C_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0C_Y07_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0B_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0B_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0B_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0B_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0B_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0B_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0B_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0B_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0B_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0B_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0A_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0A_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0B_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0B_Y07_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y07_clk_pass_through_out_right),
    .clk_out(Tile_X0B_Y07_clk_out),
    .config_config_addr(Tile_X0B_Y06_config_out_config_addr),
    .config_config_data(Tile_X0B_Y06_config_out_config_data),
    .config_out_config_addr(Tile_X0B_Y07_config_out_config_addr),
    .config_out_config_data(Tile_X0B_Y07_config_out_config_data),
    .config_out_read(Tile_X0B_Y07_config_out_read),
    .config_out_write(Tile_X0B_Y07_config_out_write),
    .config_read(Tile_X0B_Y06_config_out_read),
    .config_write(Tile_X0B_Y06_config_out_write),
    .hi(Tile_X0B_Y07_hi_unq1),
    .lo(Tile_X0B_Y07_lo_unq1),
    .read_config_data(Tile_X0B_Y07_read_config_data),
    .read_config_data_in(Tile_X0B_Y06_read_config_data),
    .reset(Tile_X0B_Y06_reset_out),
    .reset_out(Tile_X0B_Y07_reset_out),
    .stall(Tile_X0B_Y06_stall_out),
    .stall_out(Tile_X0B_Y07_stall_out),
    .tile_id(Tile_X0B_Y07_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0B_Y07_hi (
    .in(Tile_X0B_Y07_hi_unq1),
    .out(Tile_X0B_Y07_hi_out)
);
mantle_wire__typeBit8 Tile_X0B_Y07_lo (
    .in(Tile_X0B_Y07_lo_unq1),
    .out(Tile_X0B_Y07_lo_out)
);
wire [15:0] Tile_X0B_Y07_tile_id_out;
assign Tile_X0B_Y07_tile_id_out = {Tile_X0B_Y07_lo_out[7],Tile_X0B_Y07_lo_out[7:6],Tile_X0B_Y07_lo_out[6],Tile_X0B_Y07_hi_out[6],Tile_X0B_Y07_lo_out[5],Tile_X0B_Y07_hi_out[5:4],Tile_X0B_Y07_lo_out[3],Tile_X0B_Y07_lo_out[3:2],Tile_X0B_Y07_lo_out[2:1],Tile_X0B_Y07_hi_out[1],Tile_X0B_Y07_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X0B_Y07_tile_id (
    .in(Tile_X0B_Y07_tile_id_in),
    .out(Tile_X0B_Y07_tile_id_out)
);
Tile_MemCore Tile_X0B_Y08 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0C_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0C_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0B_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0B_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0B_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0B_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0B_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0B_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0B_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0B_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0B_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0B_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0A_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0A_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0B_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0B_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0C_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0C_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0B_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0B_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0B_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0B_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0B_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0B_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0B_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0B_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0B_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0B_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0A_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0A_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0B_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0B_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0C_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0C_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0B_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0B_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0B_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0B_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0B_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0B_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0B_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0B_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0B_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0B_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0A_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0A_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0B_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0B_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0C_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0C_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0B_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0B_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0B_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0B_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0B_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0B_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0B_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0B_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0B_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0B_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0A_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0A_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0B_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0B_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0C_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0C_Y08_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0B_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0B_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0B_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0B_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0B_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0B_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0B_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0B_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0B_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0B_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0A_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0A_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0B_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0B_Y08_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y08_clk_pass_through_out_right),
    .clk_out(Tile_X0B_Y08_clk_out),
    .config_config_addr(Tile_X0B_Y07_config_out_config_addr),
    .config_config_data(Tile_X0B_Y07_config_out_config_data),
    .config_out_config_addr(Tile_X0B_Y08_config_out_config_addr),
    .config_out_config_data(Tile_X0B_Y08_config_out_config_data),
    .config_out_read(Tile_X0B_Y08_config_out_read),
    .config_out_write(Tile_X0B_Y08_config_out_write),
    .config_read(Tile_X0B_Y07_config_out_read),
    .config_write(Tile_X0B_Y07_config_out_write),
    .hi(Tile_X0B_Y08_hi_unq1),
    .lo(Tile_X0B_Y08_lo_unq1),
    .read_config_data(Tile_X0B_Y08_read_config_data),
    .read_config_data_in(Tile_X0B_Y07_read_config_data),
    .reset(Tile_X0B_Y07_reset_out),
    .reset_out(Tile_X0B_Y08_reset_out),
    .stall(Tile_X0B_Y07_stall_out),
    .stall_out(Tile_X0B_Y08_stall_out),
    .tile_id(Tile_X0B_Y08_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0B_Y08_hi (
    .in(Tile_X0B_Y08_hi_unq1),
    .out(Tile_X0B_Y08_hi_out)
);
mantle_wire__typeBit8 Tile_X0B_Y08_lo (
    .in(Tile_X0B_Y08_lo_unq1),
    .out(Tile_X0B_Y08_lo_out)
);
wire [15:0] Tile_X0B_Y08_tile_id_out;
assign Tile_X0B_Y08_tile_id_out = {Tile_X0B_Y08_lo_out[7],Tile_X0B_Y08_lo_out[7:6],Tile_X0B_Y08_lo_out[6],Tile_X0B_Y08_hi_out[6],Tile_X0B_Y08_lo_out[5],Tile_X0B_Y08_hi_out[5:4],Tile_X0B_Y08_lo_out[3],Tile_X0B_Y08_lo_out[3:2],Tile_X0B_Y08_lo_out[2],Tile_X0B_Y08_hi_out[2],Tile_X0B_Y08_lo_out[1:0],Tile_X0B_Y08_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0B_Y08_tile_id (
    .in(Tile_X0B_Y08_tile_id_in),
    .out(Tile_X0B_Y08_tile_id_out)
);
Tile_MemCore Tile_X0B_Y09 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0C_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0C_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0B_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0B_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0B_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0B_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0B_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0B_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0B_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0B_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0B_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0B_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0A_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0A_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0B_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0B_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0C_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0C_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0B_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0B_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0B_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0B_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0B_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0B_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0B_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0B_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0B_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0B_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0A_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0A_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0B_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0B_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0C_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0C_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0B_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0B_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0B_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0B_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0B_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0B_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0B_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0B_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0B_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0B_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0A_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0A_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0B_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0B_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0C_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0C_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0B_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0B_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0B_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0B_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0B_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0B_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0B_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0B_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0B_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0B_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0A_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0A_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0B_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0B_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0C_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0C_Y09_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0B_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0B_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0B_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0B_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0B_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0B_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0B_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0B_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0B_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0B_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0A_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0A_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0B_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0B_Y09_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y09_clk_pass_through_out_right),
    .clk_out(Tile_X0B_Y09_clk_out),
    .config_config_addr(ConfigPipeStage_inst11_config_out_config_addr),
    .config_config_data(ConfigPipeStage_inst11_config_out_config_data),
    .config_out_config_addr(Tile_X0B_Y09_config_out_config_addr),
    .config_out_config_data(Tile_X0B_Y09_config_out_config_data),
    .config_out_read(Tile_X0B_Y09_config_out_read),
    .config_out_write(Tile_X0B_Y09_config_out_write),
    .config_read(ConfigPipeStage_inst11_config_out_read),
    .config_write(ConfigPipeStage_inst11_config_out_write),
    .hi(Tile_X0B_Y09_hi_unq1),
    .lo(Tile_X0B_Y09_lo_unq1),
    .read_config_data(Tile_X0B_Y09_read_config_data),
    .read_config_data_in(Tile_X0B_Y08_read_config_data),
    .reset(Tile_X0B_Y08_reset_out),
    .reset_out(Tile_X0B_Y09_reset_out),
    .stall(Tile_X0B_Y08_stall_out),
    .stall_out(Tile_X0B_Y09_stall_out),
    .tile_id(Tile_X0B_Y09_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0B_Y09_hi (
    .in(Tile_X0B_Y09_hi_unq1),
    .out(Tile_X0B_Y09_hi_out)
);
mantle_wire__typeBit8 Tile_X0B_Y09_lo (
    .in(Tile_X0B_Y09_lo_unq1),
    .out(Tile_X0B_Y09_lo_out)
);
wire [15:0] Tile_X0B_Y09_tile_id_out;
assign Tile_X0B_Y09_tile_id_out = {Tile_X0B_Y09_lo_out[7],Tile_X0B_Y09_lo_out[7:6],Tile_X0B_Y09_lo_out[6],Tile_X0B_Y09_hi_out[6],Tile_X0B_Y09_lo_out[5],Tile_X0B_Y09_hi_out[5:4],Tile_X0B_Y09_lo_out[3],Tile_X0B_Y09_lo_out[3:2],Tile_X0B_Y09_lo_out[2],Tile_X0B_Y09_hi_out[2],Tile_X0B_Y09_lo_out[1:0],Tile_X0B_Y09_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X0B_Y09_tile_id (
    .in(Tile_X0B_Y09_tile_id_in),
    .out(Tile_X0B_Y09_tile_id_out)
);
Tile_MemCore Tile_X0B_Y0A (
    .SB_T0_EAST_SB_IN_B1(Tile_X0C_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0C_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0B_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0B_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0B_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0B_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0B_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0B_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0B_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0B_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0B_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0B_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0A_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0A_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0B_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0B_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0C_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0C_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0B_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0B_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0B_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0B_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0B_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0B_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0B_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0B_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0B_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0B_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0A_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0A_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0B_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0B_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0C_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0C_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0B_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0B_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0B_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0B_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0B_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0B_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0B_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0B_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0B_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0B_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0A_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0A_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0B_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0B_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0C_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0C_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0B_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0B_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0B_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0B_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0B_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0B_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0B_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0B_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0B_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0B_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0A_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0A_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0B_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0B_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0C_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0C_Y0A_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0B_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0B_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0B_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0B_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0B_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0B_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0B_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0B_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0B_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0B_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0A_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0A_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0B_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0B_Y0A_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y0A_clk_pass_through_out_right),
    .clk_out(Tile_X0B_Y0A_clk_out),
    .config_config_addr(Tile_X0B_Y09_config_out_config_addr),
    .config_config_data(Tile_X0B_Y09_config_out_config_data),
    .config_out_config_addr(Tile_X0B_Y0A_config_out_config_addr),
    .config_out_config_data(Tile_X0B_Y0A_config_out_config_data),
    .config_out_read(Tile_X0B_Y0A_config_out_read),
    .config_out_write(Tile_X0B_Y0A_config_out_write),
    .config_read(Tile_X0B_Y09_config_out_read),
    .config_write(Tile_X0B_Y09_config_out_write),
    .hi(Tile_X0B_Y0A_hi_unq1),
    .lo(Tile_X0B_Y0A_lo_unq1),
    .read_config_data(Tile_X0B_Y0A_read_config_data),
    .read_config_data_in(Tile_X0B_Y09_read_config_data),
    .reset(Tile_X0B_Y09_reset_out),
    .reset_out(Tile_X0B_Y0A_reset_out),
    .stall(Tile_X0B_Y09_stall_out),
    .stall_out(Tile_X0B_Y0A_stall_out),
    .tile_id(Tile_X0B_Y0A_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0B_Y0A_hi (
    .in(Tile_X0B_Y0A_hi_unq1),
    .out(Tile_X0B_Y0A_hi_out)
);
mantle_wire__typeBit8 Tile_X0B_Y0A_lo (
    .in(Tile_X0B_Y0A_lo_unq1),
    .out(Tile_X0B_Y0A_lo_out)
);
wire [15:0] Tile_X0B_Y0A_tile_id_out;
assign Tile_X0B_Y0A_tile_id_out = {Tile_X0B_Y0A_lo_out[7],Tile_X0B_Y0A_lo_out[7:6],Tile_X0B_Y0A_lo_out[6],Tile_X0B_Y0A_hi_out[6],Tile_X0B_Y0A_lo_out[5],Tile_X0B_Y0A_hi_out[5:4],Tile_X0B_Y0A_lo_out[3],Tile_X0B_Y0A_lo_out[3:2],Tile_X0B_Y0A_lo_out[2],Tile_X0B_Y0A_hi_out[2],Tile_X0B_Y0A_lo_out[1],Tile_X0B_Y0A_hi_out[1],Tile_X0B_Y0A_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0B_Y0A_tile_id (
    .in(Tile_X0B_Y0A_tile_id_in),
    .out(Tile_X0B_Y0A_tile_id_out)
);
Tile_MemCore Tile_X0B_Y0B (
    .SB_T0_EAST_SB_IN_B1(Tile_X0C_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0C_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0B_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0B_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0B_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0B_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0B_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0B_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0B_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0B_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0B_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0B_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0A_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0A_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0B_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0B_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0C_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0C_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0B_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0B_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0B_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0B_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0B_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0B_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0B_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0B_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0B_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0B_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0A_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0A_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0B_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0B_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0C_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0C_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0B_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0B_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0B_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0B_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0B_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0B_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0B_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0B_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0B_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0B_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0A_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0A_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0B_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0B_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0C_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0C_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0B_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0B_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0B_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0B_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0B_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0B_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0B_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0B_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0B_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0B_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0A_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0A_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0B_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0B_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0C_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0C_Y0B_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0B_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0B_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0B_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0B_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0B_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0B_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0B_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0B_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0B_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0B_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0A_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0A_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0B_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0B_Y0B_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y0B_clk_pass_through_out_right),
    .clk_out(Tile_X0B_Y0B_clk_out),
    .config_config_addr(Tile_X0B_Y0A_config_out_config_addr),
    .config_config_data(Tile_X0B_Y0A_config_out_config_data),
    .config_out_config_addr(Tile_X0B_Y0B_config_out_config_addr),
    .config_out_config_data(Tile_X0B_Y0B_config_out_config_data),
    .config_out_read(Tile_X0B_Y0B_config_out_read),
    .config_out_write(Tile_X0B_Y0B_config_out_write),
    .config_read(Tile_X0B_Y0A_config_out_read),
    .config_write(Tile_X0B_Y0A_config_out_write),
    .hi(Tile_X0B_Y0B_hi_unq1),
    .lo(Tile_X0B_Y0B_lo_unq1),
    .read_config_data(Tile_X0B_Y0B_read_config_data),
    .read_config_data_in(Tile_X0B_Y0A_read_config_data),
    .reset(Tile_X0B_Y0A_reset_out),
    .reset_out(Tile_X0B_Y0B_reset_out),
    .stall(Tile_X0B_Y0A_stall_out),
    .stall_out(Tile_X0B_Y0B_stall_out),
    .tile_id(Tile_X0B_Y0B_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0B_Y0B_hi (
    .in(Tile_X0B_Y0B_hi_unq1),
    .out(Tile_X0B_Y0B_hi_out)
);
mantle_wire__typeBit8 Tile_X0B_Y0B_lo (
    .in(Tile_X0B_Y0B_lo_unq1),
    .out(Tile_X0B_Y0B_lo_out)
);
wire [15:0] Tile_X0B_Y0B_tile_id_out;
assign Tile_X0B_Y0B_tile_id_out = {Tile_X0B_Y0B_lo_out[7],Tile_X0B_Y0B_lo_out[7:6],Tile_X0B_Y0B_lo_out[6],Tile_X0B_Y0B_hi_out[6],Tile_X0B_Y0B_lo_out[5],Tile_X0B_Y0B_hi_out[5:4],Tile_X0B_Y0B_lo_out[3],Tile_X0B_Y0B_lo_out[3:2],Tile_X0B_Y0B_lo_out[2],Tile_X0B_Y0B_hi_out[2],Tile_X0B_Y0B_lo_out[1],Tile_X0B_Y0B_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X0B_Y0B_tile_id (
    .in(Tile_X0B_Y0B_tile_id_in),
    .out(Tile_X0B_Y0B_tile_id_out)
);
Tile_MemCore Tile_X0B_Y0C (
    .SB_T0_EAST_SB_IN_B1(Tile_X0C_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0C_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0B_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0B_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0B_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0B_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0B_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0B_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0B_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0B_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0B_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0B_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0A_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0A_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0B_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0B_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0C_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0C_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0B_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0B_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0B_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0B_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0B_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0B_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0B_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0B_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0B_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0B_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0A_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0A_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0B_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0B_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0C_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0C_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0B_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0B_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0B_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0B_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0B_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0B_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0B_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0B_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0B_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0B_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0A_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0A_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0B_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0B_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0C_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0C_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0B_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0B_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0B_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0B_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0B_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0B_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0B_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0B_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0B_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0B_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0A_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0A_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0B_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0B_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0C_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0C_Y0C_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0B_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0B_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0B_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0B_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0B_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0B_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0B_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0B_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0B_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0B_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0A_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0A_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0B_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0B_Y0C_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y0C_clk_pass_through_out_right),
    .clk_out(Tile_X0B_Y0C_clk_out),
    .config_config_addr(Tile_X0B_Y0B_config_out_config_addr),
    .config_config_data(Tile_X0B_Y0B_config_out_config_data),
    .config_out_config_addr(Tile_X0B_Y0C_config_out_config_addr),
    .config_out_config_data(Tile_X0B_Y0C_config_out_config_data),
    .config_out_read(Tile_X0B_Y0C_config_out_read),
    .config_out_write(Tile_X0B_Y0C_config_out_write),
    .config_read(Tile_X0B_Y0B_config_out_read),
    .config_write(Tile_X0B_Y0B_config_out_write),
    .hi(Tile_X0B_Y0C_hi_unq1),
    .lo(Tile_X0B_Y0C_lo_unq1),
    .read_config_data(Tile_X0B_Y0C_read_config_data),
    .read_config_data_in(Tile_X0B_Y0B_read_config_data),
    .reset(Tile_X0B_Y0B_reset_out),
    .reset_out(Tile_X0B_Y0C_reset_out),
    .stall(Tile_X0B_Y0B_stall_out),
    .stall_out(Tile_X0B_Y0C_stall_out),
    .tile_id(Tile_X0B_Y0C_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0B_Y0C_hi (
    .in(Tile_X0B_Y0C_hi_unq1),
    .out(Tile_X0B_Y0C_hi_out)
);
mantle_wire__typeBit8 Tile_X0B_Y0C_lo (
    .in(Tile_X0B_Y0C_lo_unq1),
    .out(Tile_X0B_Y0C_lo_out)
);
wire [15:0] Tile_X0B_Y0C_tile_id_out;
assign Tile_X0B_Y0C_tile_id_out = {Tile_X0B_Y0C_lo_out[7],Tile_X0B_Y0C_lo_out[7:6],Tile_X0B_Y0C_lo_out[6],Tile_X0B_Y0C_hi_out[6],Tile_X0B_Y0C_lo_out[5],Tile_X0B_Y0C_hi_out[5:4],Tile_X0B_Y0C_lo_out[3],Tile_X0B_Y0C_lo_out[3:2],Tile_X0B_Y0C_lo_out[2],Tile_X0B_Y0C_hi_out[2:1],Tile_X0B_Y0C_lo_out[0],Tile_X0B_Y0C_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0B_Y0C_tile_id (
    .in(Tile_X0B_Y0C_tile_id_in),
    .out(Tile_X0B_Y0C_tile_id_out)
);
Tile_MemCore Tile_X0B_Y0D (
    .SB_T0_EAST_SB_IN_B1(Tile_X0C_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0C_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0B_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0B_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0B_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0B_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0B_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0B_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0B_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0B_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0B_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0B_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0A_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0A_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0B_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0B_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0C_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0C_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0B_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0B_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0B_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0B_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0B_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0B_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0B_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0B_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0B_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0B_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0A_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0A_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0B_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0B_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0C_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0C_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0B_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0B_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0B_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0B_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0B_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0B_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0B_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0B_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0B_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0B_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0A_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0A_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0B_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0B_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0C_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0C_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0B_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0B_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0B_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0B_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0B_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0B_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0B_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0B_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0B_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0B_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0A_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0A_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0B_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0B_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0C_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0C_Y0D_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0B_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0B_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0B_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0B_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0B_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0B_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0B_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0B_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0B_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0B_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0A_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0A_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0B_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0B_Y0D_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y0D_clk_pass_through_out_right),
    .clk_out(Tile_X0B_Y0D_clk_out),
    .config_config_addr(Tile_X0B_Y0C_config_out_config_addr),
    .config_config_data(Tile_X0B_Y0C_config_out_config_data),
    .config_out_config_addr(Tile_X0B_Y0D_config_out_config_addr),
    .config_out_config_data(Tile_X0B_Y0D_config_out_config_data),
    .config_out_read(Tile_X0B_Y0D_config_out_read),
    .config_out_write(Tile_X0B_Y0D_config_out_write),
    .config_read(Tile_X0B_Y0C_config_out_read),
    .config_write(Tile_X0B_Y0C_config_out_write),
    .hi(Tile_X0B_Y0D_hi_unq1),
    .lo(Tile_X0B_Y0D_lo_unq1),
    .read_config_data(Tile_X0B_Y0D_read_config_data),
    .read_config_data_in(Tile_X0B_Y0C_read_config_data),
    .reset(Tile_X0B_Y0C_reset_out),
    .reset_out(Tile_X0B_Y0D_reset_out),
    .stall(Tile_X0B_Y0C_stall_out),
    .stall_out(Tile_X0B_Y0D_stall_out),
    .tile_id(Tile_X0B_Y0D_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0B_Y0D_hi (
    .in(Tile_X0B_Y0D_hi_unq1),
    .out(Tile_X0B_Y0D_hi_out)
);
mantle_wire__typeBit8 Tile_X0B_Y0D_lo (
    .in(Tile_X0B_Y0D_lo_unq1),
    .out(Tile_X0B_Y0D_lo_out)
);
wire [15:0] Tile_X0B_Y0D_tile_id_out;
assign Tile_X0B_Y0D_tile_id_out = {Tile_X0B_Y0D_lo_out[7],Tile_X0B_Y0D_lo_out[7:6],Tile_X0B_Y0D_lo_out[6],Tile_X0B_Y0D_hi_out[6],Tile_X0B_Y0D_lo_out[5],Tile_X0B_Y0D_hi_out[5:4],Tile_X0B_Y0D_lo_out[3],Tile_X0B_Y0D_lo_out[3:2],Tile_X0B_Y0D_lo_out[2],Tile_X0B_Y0D_hi_out[2:1],Tile_X0B_Y0D_lo_out[0],Tile_X0B_Y0D_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X0B_Y0D_tile_id (
    .in(Tile_X0B_Y0D_tile_id_in),
    .out(Tile_X0B_Y0D_tile_id_out)
);
Tile_MemCore Tile_X0B_Y0E (
    .SB_T0_EAST_SB_IN_B1(Tile_X0C_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0C_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0B_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0B_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0B_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0B_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0B_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0B_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0B_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0B_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0B_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0B_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0A_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0A_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0B_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0B_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0C_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0C_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0B_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0B_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0B_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0B_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0B_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0B_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0B_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0B_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0B_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0B_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0A_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0A_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0B_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0B_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0C_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0C_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0B_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0B_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0B_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0B_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0B_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0B_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0B_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0B_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0B_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0B_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0A_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0A_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0B_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0B_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0C_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0C_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0B_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0B_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0B_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0B_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0B_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0B_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0B_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0B_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0B_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0B_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0A_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0A_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0B_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0B_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0C_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0C_Y0E_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0B_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0B_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0B_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0B_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0B_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0B_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0B_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0B_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0B_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0B_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0A_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0A_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0B_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0B_Y0E_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y0E_clk_pass_through_out_right),
    .clk_out(Tile_X0B_Y0E_clk_out),
    .config_config_addr(Tile_X0B_Y0D_config_out_config_addr),
    .config_config_data(Tile_X0B_Y0D_config_out_config_data),
    .config_out_config_addr(Tile_X0B_Y0E_config_out_config_addr),
    .config_out_config_data(Tile_X0B_Y0E_config_out_config_data),
    .config_out_read(Tile_X0B_Y0E_config_out_read),
    .config_out_write(Tile_X0B_Y0E_config_out_write),
    .config_read(Tile_X0B_Y0D_config_out_read),
    .config_write(Tile_X0B_Y0D_config_out_write),
    .hi(Tile_X0B_Y0E_hi_unq1),
    .lo(Tile_X0B_Y0E_lo_unq1),
    .read_config_data(Tile_X0B_Y0E_read_config_data),
    .read_config_data_in(Tile_X0B_Y0D_read_config_data),
    .reset(Tile_X0B_Y0D_reset_out),
    .reset_out(Tile_X0B_Y0E_reset_out),
    .stall(Tile_X0B_Y0D_stall_out),
    .stall_out(Tile_X0B_Y0E_stall_out),
    .tile_id(Tile_X0B_Y0E_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0B_Y0E_hi (
    .in(Tile_X0B_Y0E_hi_unq1),
    .out(Tile_X0B_Y0E_hi_out)
);
mantle_wire__typeBit8 Tile_X0B_Y0E_lo (
    .in(Tile_X0B_Y0E_lo_unq1),
    .out(Tile_X0B_Y0E_lo_out)
);
wire [15:0] Tile_X0B_Y0E_tile_id_out;
assign Tile_X0B_Y0E_tile_id_out = {Tile_X0B_Y0E_lo_out[7],Tile_X0B_Y0E_lo_out[7:6],Tile_X0B_Y0E_lo_out[6],Tile_X0B_Y0E_hi_out[6],Tile_X0B_Y0E_lo_out[5],Tile_X0B_Y0E_hi_out[5:4],Tile_X0B_Y0E_lo_out[3],Tile_X0B_Y0E_lo_out[3:2],Tile_X0B_Y0E_lo_out[2],Tile_X0B_Y0E_hi_out[2:1],Tile_X0B_Y0E_hi_out[1],Tile_X0B_Y0E_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0B_Y0E_tile_id (
    .in(Tile_X0B_Y0E_tile_id_in),
    .out(Tile_X0B_Y0E_tile_id_out)
);
Tile_MemCore Tile_X0B_Y0F (
    .SB_T0_EAST_SB_IN_B1(Tile_X0C_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0C_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0B_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0B_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0B_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0B_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0B_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0B_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0B_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0B_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0B_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0B_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0A_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0A_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0B_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0B_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0C_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0C_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0B_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0B_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0B_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0B_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0B_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0B_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0B_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0B_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0B_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0B_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0A_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0A_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0B_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0B_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0C_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0C_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0B_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0B_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0B_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0B_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0B_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0B_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0B_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0B_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0B_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0B_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0A_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0A_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0B_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0B_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0C_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0C_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0B_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0B_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0B_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0B_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0B_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0B_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0B_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0B_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0B_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0B_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0A_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0A_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0B_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0B_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0C_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0C_Y0F_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0B_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0B_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0B_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0B_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0B_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0B_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0B_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0B_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0B_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0B_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0A_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0A_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0B_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0B_Y0F_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y0F_clk_pass_through_out_right),
    .clk_out(Tile_X0B_Y0F_clk_out),
    .config_config_addr(Tile_X0B_Y0E_config_out_config_addr),
    .config_config_data(Tile_X0B_Y0E_config_out_config_data),
    .config_out_config_addr(Tile_X0B_Y0F_config_out_config_addr),
    .config_out_config_data(Tile_X0B_Y0F_config_out_config_data),
    .config_out_read(Tile_X0B_Y0F_config_out_read),
    .config_out_write(Tile_X0B_Y0F_config_out_write),
    .config_read(Tile_X0B_Y0E_config_out_read),
    .config_write(Tile_X0B_Y0E_config_out_write),
    .hi(Tile_X0B_Y0F_hi_unq1),
    .lo(Tile_X0B_Y0F_lo_unq1),
    .read_config_data(Tile_X0B_Y0F_read_config_data),
    .read_config_data_in(Tile_X0B_Y0E_read_config_data),
    .reset(Tile_X0B_Y0E_reset_out),
    .reset_out(Tile_X0B_Y0F_reset_out),
    .stall(Tile_X0B_Y0E_stall_out),
    .stall_out(Tile_X0B_Y0F_stall_out),
    .tile_id(Tile_X0B_Y0F_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0B_Y0F_hi (
    .in(Tile_X0B_Y0F_hi_unq1),
    .out(Tile_X0B_Y0F_hi_out)
);
mantle_wire__typeBit8 Tile_X0B_Y0F_lo (
    .in(Tile_X0B_Y0F_lo_unq1),
    .out(Tile_X0B_Y0F_lo_out)
);
wire [15:0] Tile_X0B_Y0F_tile_id_out;
assign Tile_X0B_Y0F_tile_id_out = {Tile_X0B_Y0F_lo_out[7],Tile_X0B_Y0F_lo_out[7:6],Tile_X0B_Y0F_lo_out[6],Tile_X0B_Y0F_hi_out[6],Tile_X0B_Y0F_lo_out[5],Tile_X0B_Y0F_hi_out[5:4],Tile_X0B_Y0F_lo_out[3],Tile_X0B_Y0F_lo_out[3:2],Tile_X0B_Y0F_lo_out[2],Tile_X0B_Y0F_hi_out[2:1],Tile_X0B_Y0F_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X0B_Y0F_tile_id (
    .in(Tile_X0B_Y0F_tile_id_in),
    .out(Tile_X0B_Y0F_tile_id_out)
);
Tile_MemCore Tile_X0B_Y10 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0C_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0C_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0B_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0B_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0B_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0B_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0B_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0B_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T0_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0B_Y10_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0B_Y10_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0A_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0A_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0B_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0B_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0C_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0C_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0B_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0B_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0B_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0B_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0B_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0B_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T1_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0B_Y10_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0B_Y10_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0A_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0A_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0B_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0B_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0C_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0C_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0B_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0B_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0B_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0B_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0B_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0B_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T2_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0B_Y10_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0B_Y10_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0A_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0A_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0B_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0B_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0C_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0C_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0B_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0B_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0B_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0B_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0B_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0B_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T3_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0B_Y10_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0B_Y10_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0A_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0A_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0B_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0B_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0C_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0C_Y10_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0B_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0B_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0B_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0B_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0B_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0B_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T4_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0B_Y10_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0B_Y10_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0A_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0A_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0B_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0B_Y10_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0A_Y10_clk_pass_through_out_right),
    .clk_out(Tile_X0B_Y10_clk_out),
    .config_config_addr(Tile_X0B_Y0F_config_out_config_addr),
    .config_config_data(Tile_X0B_Y0F_config_out_config_data),
    .config_out_config_addr(Tile_X0B_Y10_config_out_config_addr),
    .config_out_config_data(Tile_X0B_Y10_config_out_config_data),
    .config_out_read(Tile_X0B_Y10_config_out_read),
    .config_out_write(Tile_X0B_Y10_config_out_write),
    .config_read(Tile_X0B_Y0F_config_out_read),
    .config_write(Tile_X0B_Y0F_config_out_write),
    .hi(Tile_X0B_Y10_hi_unq1),
    .lo(Tile_X0B_Y10_lo_unq1),
    .read_config_data(Tile_X0B_Y10_read_config_data),
    .read_config_data_in(Tile_X0B_Y0F_read_config_data),
    .reset(Tile_X0B_Y0F_reset_out),
    .reset_out(Tile_X0B_Y10_reset_out),
    .stall(Tile_X0B_Y0F_stall_out),
    .stall_out(Tile_X0B_Y10_stall_out),
    .tile_id(Tile_X0B_Y10_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0B_Y10_hi (
    .in(Tile_X0B_Y10_hi_unq1),
    .out(Tile_X0B_Y10_hi_out)
);
mantle_wire__typeBit8 Tile_X0B_Y10_lo (
    .in(Tile_X0B_Y10_lo_unq1),
    .out(Tile_X0B_Y10_lo_out)
);
wire [15:0] Tile_X0B_Y10_tile_id_out;
assign Tile_X0B_Y10_tile_id_out = {Tile_X0B_Y10_lo_out[7],Tile_X0B_Y10_lo_out[7:6],Tile_X0B_Y10_lo_out[6],Tile_X0B_Y10_hi_out[6],Tile_X0B_Y10_lo_out[5],Tile_X0B_Y10_hi_out[5:4],Tile_X0B_Y10_lo_out[3],Tile_X0B_Y10_lo_out[3:2],Tile_X0B_Y10_hi_out[2],Tile_X0B_Y10_lo_out[1],Tile_X0B_Y10_lo_out[1:0],Tile_X0B_Y10_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0B_Y10_tile_id (
    .in(Tile_X0B_Y10_tile_id_in),
    .out(Tile_X0B_Y10_tile_id_out)
);
wire [15:0] Tile_X0C_Y00_tile_id;
assign Tile_X0C_Y00_tile_id = {Tile_X0C_Y00_lo[7],Tile_X0C_Y00_lo[7:6],Tile_X0C_Y00_lo[6],Tile_X0C_Y00_hi[6:5],Tile_X0C_Y00_lo[4],Tile_X0C_Y00_lo[4:3],Tile_X0C_Y00_lo[3:2],Tile_X0C_Y00_lo[2:1],Tile_X0C_Y00_lo[1:0],Tile_X0C_Y00_lo[0]};
Tile_io_core Tile_X0C_Y00 (
    .tile_id(Tile_X0C_Y00_tile_id),
    .glb2io_1(glb2io_1_X0C_Y00),
    .f2io_1(Tile_X0C_Y01_SB_T0_NORTH_SB_OUT_B1),
    .io2glb_1(Tile_X0C_Y00_io2glb_1),
    .io2f_1(Tile_X0C_Y00_io2f_1),
    .glb2io_16(glb2io_16_X0C_Y00),
    .f2io_16(Tile_X0C_Y01_SB_T0_NORTH_SB_OUT_B16),
    .io2glb_16(Tile_X0C_Y00_io2glb_16),
    .io2f_16(Tile_X0C_Y00_io2f_16),
    .hi(Tile_X0C_Y00_hi),
    .lo(Tile_X0C_Y00_lo)
);
Tile_PE Tile_X0C_Y01 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0D_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0D_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0C_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0C_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0C_Y00_io2f_1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0C_Y00_io2f_16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0C_Y01_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0C_Y01_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0C_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0C_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0C_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0C_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0B_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0B_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0C_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0C_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0D_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0D_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0C_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0C_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0C_Y00_io2f_1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0C_Y00_io2f_16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0C_Y01_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0C_Y01_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0C_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0C_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0C_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0C_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0B_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0B_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0C_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0C_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0D_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0D_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0C_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0C_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0C_Y00_io2f_1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0C_Y00_io2f_16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0C_Y01_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0C_Y01_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0C_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0C_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0C_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0C_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0B_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0B_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0C_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0C_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0D_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0D_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0C_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0C_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0C_Y00_io2f_1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0C_Y00_io2f_16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0C_Y01_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0C_Y01_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0C_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0C_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0C_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0C_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0B_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0B_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0C_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0C_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0D_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0D_Y01_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0C_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0C_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0C_Y00_io2f_1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0C_Y00_io2f_16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0C_Y01_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0C_Y01_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0C_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0C_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0C_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0C_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0B_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0B_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0C_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0C_Y01_SB_T4_WEST_SB_OUT_B16),
    .clk(clk),
    .clk_out(Tile_X0C_Y01_clk_out),
    .clk_pass_through(clk),
    .clk_pass_through_out_bot(Tile_X0C_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0C_Y01_clk_pass_through_out_right),
    .config_config_addr(config_12_config_addr),
    .config_config_data(config_12_config_data),
    .config_out_config_addr(Tile_X0C_Y01_config_out_config_addr),
    .config_out_config_data(Tile_X0C_Y01_config_out_config_data),
    .config_out_read(Tile_X0C_Y01_config_out_read),
    .config_out_write(Tile_X0C_Y01_config_out_write),
    .config_read(config_12_read),
    .config_write(config_12_write),
    .hi(Tile_X0C_Y01_hi_unq1),
    .lo(Tile_X0C_Y01_lo_unq1),
    .read_config_data(Tile_X0C_Y01_read_config_data),
    .read_config_data_in(const_0_32_out),
    .reset(reset),
    .reset_out(Tile_X0C_Y01_reset_out),
    .stall(stall[12]),
    .stall_out(Tile_X0C_Y01_stall_out),
    .tile_id(Tile_X0C_Y01_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0C_Y01_hi (
    .in(Tile_X0C_Y01_hi_unq1),
    .out(Tile_X0C_Y01_hi_out)
);
mantle_wire__typeBit8 Tile_X0C_Y01_lo (
    .in(Tile_X0C_Y01_lo_unq1),
    .out(Tile_X0C_Y01_lo_out)
);
wire [15:0] Tile_X0C_Y01_tile_id_out;
assign Tile_X0C_Y01_tile_id_out = {Tile_X0C_Y01_lo_out[7],Tile_X0C_Y01_lo_out[7:6],Tile_X0C_Y01_lo_out[6],Tile_X0C_Y01_hi_out[6:5],Tile_X0C_Y01_lo_out[4],Tile_X0C_Y01_lo_out[4:3],Tile_X0C_Y01_lo_out[3:2],Tile_X0C_Y01_lo_out[2:1],Tile_X0C_Y01_lo_out[1:0],Tile_X0C_Y01_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X0C_Y01_tile_id (
    .in(Tile_X0C_Y01_tile_id_in),
    .out(Tile_X0C_Y01_tile_id_out)
);
Tile_PE Tile_X0C_Y02 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0D_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0D_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0C_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0C_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0C_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0C_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0C_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0C_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0C_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0C_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0C_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0C_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0B_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0B_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0C_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0C_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0D_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0D_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0C_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0C_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0C_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0C_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0C_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0C_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0C_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0C_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0C_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0C_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0B_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0B_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0C_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0C_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0D_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0D_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0C_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0C_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0C_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0C_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0C_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0C_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0C_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0C_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0C_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0C_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0B_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0B_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0C_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0C_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0D_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0D_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0C_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0C_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0C_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0C_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0C_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0C_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0C_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0C_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0C_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0C_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0B_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0B_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0C_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0C_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0D_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0D_Y02_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0C_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0C_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0C_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0C_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0C_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0C_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0C_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0C_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0C_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0C_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0B_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0B_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0C_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0C_Y02_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0C_Y01_clk_out),
    .clk_out(Tile_X0C_Y02_clk_out),
    .clk_pass_through(Tile_X0C_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0C_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0C_Y02_clk_pass_through_out_right),
    .config_config_addr(Tile_X0C_Y01_config_out_config_addr),
    .config_config_data(Tile_X0C_Y01_config_out_config_data),
    .config_out_config_addr(Tile_X0C_Y02_config_out_config_addr),
    .config_out_config_data(Tile_X0C_Y02_config_out_config_data),
    .config_out_read(Tile_X0C_Y02_config_out_read),
    .config_out_write(Tile_X0C_Y02_config_out_write),
    .config_read(Tile_X0C_Y01_config_out_read),
    .config_write(Tile_X0C_Y01_config_out_write),
    .hi(Tile_X0C_Y02_hi_unq1),
    .lo(Tile_X0C_Y02_lo_unq1),
    .read_config_data(Tile_X0C_Y02_read_config_data),
    .read_config_data_in(Tile_X0C_Y01_read_config_data),
    .reset(Tile_X0C_Y01_reset_out),
    .reset_out(Tile_X0C_Y02_reset_out),
    .stall(Tile_X0C_Y01_stall_out),
    .stall_out(Tile_X0C_Y02_stall_out),
    .tile_id(Tile_X0C_Y02_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0C_Y02_hi (
    .in(Tile_X0C_Y02_hi_unq1),
    .out(Tile_X0C_Y02_hi_out)
);
mantle_wire__typeBit8 Tile_X0C_Y02_lo (
    .in(Tile_X0C_Y02_lo_unq1),
    .out(Tile_X0C_Y02_lo_out)
);
wire [15:0] Tile_X0C_Y02_tile_id_out;
assign Tile_X0C_Y02_tile_id_out = {Tile_X0C_Y02_lo_out[7],Tile_X0C_Y02_lo_out[7:6],Tile_X0C_Y02_lo_out[6],Tile_X0C_Y02_hi_out[6:5],Tile_X0C_Y02_lo_out[4],Tile_X0C_Y02_lo_out[4:3],Tile_X0C_Y02_lo_out[3:2],Tile_X0C_Y02_lo_out[2:1],Tile_X0C_Y02_lo_out[1],Tile_X0C_Y02_hi_out[1],Tile_X0C_Y02_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0C_Y02_tile_id (
    .in(Tile_X0C_Y02_tile_id_in),
    .out(Tile_X0C_Y02_tile_id_out)
);
Tile_PE Tile_X0C_Y03 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0D_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0D_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0C_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0C_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0C_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0C_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0C_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0C_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0C_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0C_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0C_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0C_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0B_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0B_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0C_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0C_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0D_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0D_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0C_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0C_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0C_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0C_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0C_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0C_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0C_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0C_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0C_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0C_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0B_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0B_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0C_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0C_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0D_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0D_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0C_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0C_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0C_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0C_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0C_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0C_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0C_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0C_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0C_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0C_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0B_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0B_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0C_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0C_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0D_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0D_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0C_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0C_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0C_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0C_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0C_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0C_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0C_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0C_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0C_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0C_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0B_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0B_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0C_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0C_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0D_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0D_Y03_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0C_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0C_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0C_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0C_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0C_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0C_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0C_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0C_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0C_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0C_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0B_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0B_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0C_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0C_Y03_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0C_Y02_clk_out),
    .clk_out(Tile_X0C_Y03_clk_out),
    .clk_pass_through(Tile_X0C_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0C_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0C_Y03_clk_pass_through_out_right),
    .config_config_addr(Tile_X0C_Y02_config_out_config_addr),
    .config_config_data(Tile_X0C_Y02_config_out_config_data),
    .config_out_config_addr(Tile_X0C_Y03_config_out_config_addr),
    .config_out_config_data(Tile_X0C_Y03_config_out_config_data),
    .config_out_read(Tile_X0C_Y03_config_out_read),
    .config_out_write(Tile_X0C_Y03_config_out_write),
    .config_read(Tile_X0C_Y02_config_out_read),
    .config_write(Tile_X0C_Y02_config_out_write),
    .hi(Tile_X0C_Y03_hi_unq1),
    .lo(Tile_X0C_Y03_lo_unq1),
    .read_config_data(Tile_X0C_Y03_read_config_data),
    .read_config_data_in(Tile_X0C_Y02_read_config_data),
    .reset(Tile_X0C_Y02_reset_out),
    .reset_out(Tile_X0C_Y03_reset_out),
    .stall(Tile_X0C_Y02_stall_out),
    .stall_out(Tile_X0C_Y03_stall_out),
    .tile_id(Tile_X0C_Y03_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0C_Y03_hi (
    .in(Tile_X0C_Y03_hi_unq1),
    .out(Tile_X0C_Y03_hi_out)
);
mantle_wire__typeBit8 Tile_X0C_Y03_lo (
    .in(Tile_X0C_Y03_lo_unq1),
    .out(Tile_X0C_Y03_lo_out)
);
wire [15:0] Tile_X0C_Y03_tile_id_out;
assign Tile_X0C_Y03_tile_id_out = {Tile_X0C_Y03_lo_out[7],Tile_X0C_Y03_lo_out[7:6],Tile_X0C_Y03_lo_out[6],Tile_X0C_Y03_hi_out[6:5],Tile_X0C_Y03_lo_out[4],Tile_X0C_Y03_lo_out[4:3],Tile_X0C_Y03_lo_out[3:2],Tile_X0C_Y03_lo_out[2:1],Tile_X0C_Y03_lo_out[1],Tile_X0C_Y03_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X0C_Y03_tile_id (
    .in(Tile_X0C_Y03_tile_id_in),
    .out(Tile_X0C_Y03_tile_id_out)
);
Tile_PE Tile_X0C_Y04 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0D_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0D_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0C_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0C_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0C_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0C_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0C_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0C_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0C_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0C_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0C_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0C_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0B_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0B_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0C_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0C_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0D_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0D_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0C_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0C_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0C_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0C_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0C_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0C_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0C_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0C_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0C_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0C_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0B_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0B_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0C_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0C_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0D_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0D_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0C_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0C_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0C_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0C_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0C_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0C_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0C_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0C_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0C_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0C_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0B_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0B_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0C_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0C_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0D_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0D_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0C_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0C_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0C_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0C_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0C_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0C_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0C_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0C_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0C_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0C_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0B_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0B_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0C_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0C_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0D_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0D_Y04_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0C_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0C_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0C_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0C_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0C_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0C_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0C_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0C_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0C_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0C_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0B_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0B_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0C_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0C_Y04_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0C_Y03_clk_out),
    .clk_out(Tile_X0C_Y04_clk_out),
    .clk_pass_through(Tile_X0C_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0C_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0C_Y04_clk_pass_through_out_right),
    .config_config_addr(Tile_X0C_Y03_config_out_config_addr),
    .config_config_data(Tile_X0C_Y03_config_out_config_data),
    .config_out_config_addr(Tile_X0C_Y04_config_out_config_addr),
    .config_out_config_data(Tile_X0C_Y04_config_out_config_data),
    .config_out_read(Tile_X0C_Y04_config_out_read),
    .config_out_write(Tile_X0C_Y04_config_out_write),
    .config_read(Tile_X0C_Y03_config_out_read),
    .config_write(Tile_X0C_Y03_config_out_write),
    .hi(Tile_X0C_Y04_hi_unq1),
    .lo(Tile_X0C_Y04_lo_unq1),
    .read_config_data(Tile_X0C_Y04_read_config_data),
    .read_config_data_in(Tile_X0C_Y03_read_config_data),
    .reset(Tile_X0C_Y03_reset_out),
    .reset_out(Tile_X0C_Y04_reset_out),
    .stall(Tile_X0C_Y03_stall_out),
    .stall_out(Tile_X0C_Y04_stall_out),
    .tile_id(Tile_X0C_Y04_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0C_Y04_hi (
    .in(Tile_X0C_Y04_hi_unq1),
    .out(Tile_X0C_Y04_hi_out)
);
mantle_wire__typeBit8 Tile_X0C_Y04_lo (
    .in(Tile_X0C_Y04_lo_unq1),
    .out(Tile_X0C_Y04_lo_out)
);
wire [15:0] Tile_X0C_Y04_tile_id_out;
assign Tile_X0C_Y04_tile_id_out = {Tile_X0C_Y04_lo_out[7],Tile_X0C_Y04_lo_out[7:6],Tile_X0C_Y04_lo_out[6],Tile_X0C_Y04_hi_out[6:5],Tile_X0C_Y04_lo_out[4],Tile_X0C_Y04_lo_out[4:3],Tile_X0C_Y04_lo_out[3:2],Tile_X0C_Y04_lo_out[2:1],Tile_X0C_Y04_hi_out[1],Tile_X0C_Y04_lo_out[0],Tile_X0C_Y04_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0C_Y04_tile_id (
    .in(Tile_X0C_Y04_tile_id_in),
    .out(Tile_X0C_Y04_tile_id_out)
);
Tile_PE Tile_X0C_Y05 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0D_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0D_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0C_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0C_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0C_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0C_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0C_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0C_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0C_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0C_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0C_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0C_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0B_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0B_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0C_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0C_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0D_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0D_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0C_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0C_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0C_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0C_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0C_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0C_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0C_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0C_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0C_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0C_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0B_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0B_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0C_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0C_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0D_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0D_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0C_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0C_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0C_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0C_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0C_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0C_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0C_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0C_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0C_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0C_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0B_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0B_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0C_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0C_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0D_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0D_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0C_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0C_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0C_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0C_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0C_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0C_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0C_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0C_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0C_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0C_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0B_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0B_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0C_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0C_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0D_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0D_Y05_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0C_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0C_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0C_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0C_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0C_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0C_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0C_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0C_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0C_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0C_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0B_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0B_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0C_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0C_Y05_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0C_Y04_clk_out),
    .clk_out(Tile_X0C_Y05_clk_out),
    .clk_pass_through(Tile_X0C_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0C_Y05_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0C_Y05_clk_pass_through_out_right),
    .config_config_addr(Tile_X0C_Y04_config_out_config_addr),
    .config_config_data(Tile_X0C_Y04_config_out_config_data),
    .config_out_config_addr(Tile_X0C_Y05_config_out_config_addr),
    .config_out_config_data(Tile_X0C_Y05_config_out_config_data),
    .config_out_read(Tile_X0C_Y05_config_out_read),
    .config_out_write(Tile_X0C_Y05_config_out_write),
    .config_read(Tile_X0C_Y04_config_out_read),
    .config_write(Tile_X0C_Y04_config_out_write),
    .hi(Tile_X0C_Y05_hi_unq1),
    .lo(Tile_X0C_Y05_lo_unq1),
    .read_config_data(Tile_X0C_Y05_read_config_data),
    .read_config_data_in(Tile_X0C_Y04_read_config_data),
    .reset(Tile_X0C_Y04_reset_out),
    .reset_out(Tile_X0C_Y05_reset_out),
    .stall(Tile_X0C_Y04_stall_out),
    .stall_out(Tile_X0C_Y05_stall_out),
    .tile_id(Tile_X0C_Y05_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0C_Y05_hi (
    .in(Tile_X0C_Y05_hi_unq1),
    .out(Tile_X0C_Y05_hi_out)
);
mantle_wire__typeBit8 Tile_X0C_Y05_lo (
    .in(Tile_X0C_Y05_lo_unq1),
    .out(Tile_X0C_Y05_lo_out)
);
wire [15:0] Tile_X0C_Y05_tile_id_out;
assign Tile_X0C_Y05_tile_id_out = {Tile_X0C_Y05_lo_out[7],Tile_X0C_Y05_lo_out[7:6],Tile_X0C_Y05_lo_out[6],Tile_X0C_Y05_hi_out[6:5],Tile_X0C_Y05_lo_out[4],Tile_X0C_Y05_lo_out[4:3],Tile_X0C_Y05_lo_out[3:2],Tile_X0C_Y05_lo_out[2:1],Tile_X0C_Y05_hi_out[1],Tile_X0C_Y05_lo_out[0],Tile_X0C_Y05_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X0C_Y05_tile_id (
    .in(Tile_X0C_Y05_tile_id_in),
    .out(Tile_X0C_Y05_tile_id_out)
);
Tile_PE Tile_X0C_Y06 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0D_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0D_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0C_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0C_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0C_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0C_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0C_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0C_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0C_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0C_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0C_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0C_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0B_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0B_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0C_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0C_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0D_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0D_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0C_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0C_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0C_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0C_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0C_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0C_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0C_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0C_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0C_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0C_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0B_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0B_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0C_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0C_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0D_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0D_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0C_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0C_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0C_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0C_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0C_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0C_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0C_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0C_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0C_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0C_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0B_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0B_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0C_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0C_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0D_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0D_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0C_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0C_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0C_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0C_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0C_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0C_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0C_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0C_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0C_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0C_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0B_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0B_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0C_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0C_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0D_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0D_Y06_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0C_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0C_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0C_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0C_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0C_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0C_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0C_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0C_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0C_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0C_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0B_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0B_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0C_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0C_Y06_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0C_Y05_clk_out),
    .clk_out(Tile_X0C_Y06_clk_out),
    .clk_pass_through(Tile_X0C_Y05_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0C_Y06_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0C_Y06_clk_pass_through_out_right),
    .config_config_addr(Tile_X0C_Y05_config_out_config_addr),
    .config_config_data(Tile_X0C_Y05_config_out_config_data),
    .config_out_config_addr(Tile_X0C_Y06_config_out_config_addr),
    .config_out_config_data(Tile_X0C_Y06_config_out_config_data),
    .config_out_read(Tile_X0C_Y06_config_out_read),
    .config_out_write(Tile_X0C_Y06_config_out_write),
    .config_read(Tile_X0C_Y05_config_out_read),
    .config_write(Tile_X0C_Y05_config_out_write),
    .hi(Tile_X0C_Y06_hi_unq1),
    .lo(Tile_X0C_Y06_lo_unq1),
    .read_config_data(Tile_X0C_Y06_read_config_data),
    .read_config_data_in(Tile_X0C_Y05_read_config_data),
    .reset(Tile_X0C_Y05_reset_out),
    .reset_out(Tile_X0C_Y06_reset_out),
    .stall(Tile_X0C_Y05_stall_out),
    .stall_out(Tile_X0C_Y06_stall_out),
    .tile_id(Tile_X0C_Y06_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0C_Y06_hi (
    .in(Tile_X0C_Y06_hi_unq1),
    .out(Tile_X0C_Y06_hi_out)
);
mantle_wire__typeBit8 Tile_X0C_Y06_lo (
    .in(Tile_X0C_Y06_lo_unq1),
    .out(Tile_X0C_Y06_lo_out)
);
wire [15:0] Tile_X0C_Y06_tile_id_out;
assign Tile_X0C_Y06_tile_id_out = {Tile_X0C_Y06_lo_out[7],Tile_X0C_Y06_lo_out[7:6],Tile_X0C_Y06_lo_out[6],Tile_X0C_Y06_hi_out[6:5],Tile_X0C_Y06_lo_out[4],Tile_X0C_Y06_lo_out[4:3],Tile_X0C_Y06_lo_out[3:2],Tile_X0C_Y06_lo_out[2:1],Tile_X0C_Y06_hi_out[1],Tile_X0C_Y06_hi_out[1],Tile_X0C_Y06_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0C_Y06_tile_id (
    .in(Tile_X0C_Y06_tile_id_in),
    .out(Tile_X0C_Y06_tile_id_out)
);
Tile_PE Tile_X0C_Y07 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0D_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0D_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0C_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0C_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0C_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0C_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0C_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0C_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0C_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0C_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0C_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0C_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0B_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0B_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0C_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0C_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0D_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0D_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0C_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0C_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0C_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0C_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0C_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0C_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0C_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0C_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0C_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0C_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0B_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0B_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0C_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0C_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0D_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0D_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0C_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0C_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0C_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0C_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0C_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0C_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0C_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0C_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0C_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0C_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0B_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0B_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0C_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0C_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0D_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0D_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0C_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0C_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0C_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0C_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0C_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0C_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0C_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0C_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0C_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0C_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0B_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0B_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0C_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0C_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0D_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0D_Y07_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0C_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0C_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0C_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0C_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0C_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0C_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0C_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0C_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0C_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0C_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0B_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0B_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0C_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0C_Y07_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0C_Y06_clk_out),
    .clk_out(Tile_X0C_Y07_clk_out),
    .clk_pass_through(Tile_X0C_Y06_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0C_Y07_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0C_Y07_clk_pass_through_out_right),
    .config_config_addr(Tile_X0C_Y06_config_out_config_addr),
    .config_config_data(Tile_X0C_Y06_config_out_config_data),
    .config_out_config_addr(Tile_X0C_Y07_config_out_config_addr),
    .config_out_config_data(Tile_X0C_Y07_config_out_config_data),
    .config_out_read(Tile_X0C_Y07_config_out_read),
    .config_out_write(Tile_X0C_Y07_config_out_write),
    .config_read(Tile_X0C_Y06_config_out_read),
    .config_write(Tile_X0C_Y06_config_out_write),
    .hi(Tile_X0C_Y07_hi_unq1),
    .lo(Tile_X0C_Y07_lo_unq1),
    .read_config_data(Tile_X0C_Y07_read_config_data),
    .read_config_data_in(Tile_X0C_Y06_read_config_data),
    .reset(Tile_X0C_Y06_reset_out),
    .reset_out(Tile_X0C_Y07_reset_out),
    .stall(Tile_X0C_Y06_stall_out),
    .stall_out(Tile_X0C_Y07_stall_out),
    .tile_id(Tile_X0C_Y07_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0C_Y07_hi (
    .in(Tile_X0C_Y07_hi_unq1),
    .out(Tile_X0C_Y07_hi_out)
);
mantle_wire__typeBit8 Tile_X0C_Y07_lo (
    .in(Tile_X0C_Y07_lo_unq1),
    .out(Tile_X0C_Y07_lo_out)
);
wire [15:0] Tile_X0C_Y07_tile_id_out;
assign Tile_X0C_Y07_tile_id_out = {Tile_X0C_Y07_lo_out[7],Tile_X0C_Y07_lo_out[7:6],Tile_X0C_Y07_lo_out[6],Tile_X0C_Y07_hi_out[6:5],Tile_X0C_Y07_lo_out[4],Tile_X0C_Y07_lo_out[4:3],Tile_X0C_Y07_lo_out[3:2],Tile_X0C_Y07_lo_out[2:1],Tile_X0C_Y07_hi_out[1],Tile_X0C_Y07_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X0C_Y07_tile_id (
    .in(Tile_X0C_Y07_tile_id_in),
    .out(Tile_X0C_Y07_tile_id_out)
);
Tile_PE Tile_X0C_Y08 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0D_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0D_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0C_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0C_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0C_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0C_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0C_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0C_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0C_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0C_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0C_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0C_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0B_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0B_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0C_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0C_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0D_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0D_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0C_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0C_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0C_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0C_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0C_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0C_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0C_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0C_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0C_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0C_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0B_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0B_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0C_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0C_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0D_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0D_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0C_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0C_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0C_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0C_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0C_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0C_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0C_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0C_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0C_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0C_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0B_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0B_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0C_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0C_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0D_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0D_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0C_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0C_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0C_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0C_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0C_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0C_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0C_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0C_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0C_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0C_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0B_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0B_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0C_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0C_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0D_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0D_Y08_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0C_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0C_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0C_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0C_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0C_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0C_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0C_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0C_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0C_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0C_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0B_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0B_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0C_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0C_Y08_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0C_Y07_clk_out),
    .clk_out(Tile_X0C_Y08_clk_out),
    .clk_pass_through(Tile_X0C_Y07_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0C_Y08_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0C_Y08_clk_pass_through_out_right),
    .config_config_addr(Tile_X0C_Y07_config_out_config_addr),
    .config_config_data(Tile_X0C_Y07_config_out_config_data),
    .config_out_config_addr(Tile_X0C_Y08_config_out_config_addr),
    .config_out_config_data(Tile_X0C_Y08_config_out_config_data),
    .config_out_read(Tile_X0C_Y08_config_out_read),
    .config_out_write(Tile_X0C_Y08_config_out_write),
    .config_read(Tile_X0C_Y07_config_out_read),
    .config_write(Tile_X0C_Y07_config_out_write),
    .hi(Tile_X0C_Y08_hi_unq1),
    .lo(Tile_X0C_Y08_lo_unq1),
    .read_config_data(Tile_X0C_Y08_read_config_data),
    .read_config_data_in(Tile_X0C_Y07_read_config_data),
    .reset(Tile_X0C_Y07_reset_out),
    .reset_out(Tile_X0C_Y08_reset_out),
    .stall(Tile_X0C_Y07_stall_out),
    .stall_out(Tile_X0C_Y08_stall_out),
    .tile_id(Tile_X0C_Y08_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0C_Y08_hi (
    .in(Tile_X0C_Y08_hi_unq1),
    .out(Tile_X0C_Y08_hi_out)
);
mantle_wire__typeBit8 Tile_X0C_Y08_lo (
    .in(Tile_X0C_Y08_lo_unq1),
    .out(Tile_X0C_Y08_lo_out)
);
wire [15:0] Tile_X0C_Y08_tile_id_out;
assign Tile_X0C_Y08_tile_id_out = {Tile_X0C_Y08_lo_out[7],Tile_X0C_Y08_lo_out[7:6],Tile_X0C_Y08_lo_out[6],Tile_X0C_Y08_hi_out[6:5],Tile_X0C_Y08_lo_out[4],Tile_X0C_Y08_lo_out[4:3],Tile_X0C_Y08_lo_out[3:2],Tile_X0C_Y08_lo_out[2],Tile_X0C_Y08_hi_out[2],Tile_X0C_Y08_lo_out[1:0],Tile_X0C_Y08_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0C_Y08_tile_id (
    .in(Tile_X0C_Y08_tile_id_in),
    .out(Tile_X0C_Y08_tile_id_out)
);
Tile_PE Tile_X0C_Y09 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0D_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0D_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0C_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0C_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0C_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0C_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0C_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0C_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0C_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0C_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0C_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0C_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0B_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0B_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0C_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0C_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0D_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0D_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0C_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0C_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0C_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0C_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0C_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0C_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0C_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0C_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0C_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0C_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0B_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0B_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0C_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0C_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0D_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0D_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0C_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0C_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0C_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0C_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0C_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0C_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0C_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0C_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0C_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0C_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0B_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0B_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0C_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0C_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0D_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0D_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0C_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0C_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0C_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0C_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0C_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0C_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0C_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0C_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0C_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0C_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0B_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0B_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0C_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0C_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0D_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0D_Y09_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0C_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0C_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0C_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0C_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0C_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0C_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0C_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0C_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0C_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0C_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0B_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0B_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0C_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0C_Y09_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0C_Y08_clk_out),
    .clk_out(Tile_X0C_Y09_clk_out),
    .clk_pass_through(Tile_X0C_Y08_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0C_Y09_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0C_Y09_clk_pass_through_out_right),
    .config_config_addr(ConfigPipeStage_inst12_config_out_config_addr),
    .config_config_data(ConfigPipeStage_inst12_config_out_config_data),
    .config_out_config_addr(Tile_X0C_Y09_config_out_config_addr),
    .config_out_config_data(Tile_X0C_Y09_config_out_config_data),
    .config_out_read(Tile_X0C_Y09_config_out_read),
    .config_out_write(Tile_X0C_Y09_config_out_write),
    .config_read(ConfigPipeStage_inst12_config_out_read),
    .config_write(ConfigPipeStage_inst12_config_out_write),
    .hi(Tile_X0C_Y09_hi_unq1),
    .lo(Tile_X0C_Y09_lo_unq1),
    .read_config_data(Tile_X0C_Y09_read_config_data),
    .read_config_data_in(Tile_X0C_Y08_read_config_data),
    .reset(Tile_X0C_Y08_reset_out),
    .reset_out(Tile_X0C_Y09_reset_out),
    .stall(Tile_X0C_Y08_stall_out),
    .stall_out(Tile_X0C_Y09_stall_out),
    .tile_id(Tile_X0C_Y09_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0C_Y09_hi (
    .in(Tile_X0C_Y09_hi_unq1),
    .out(Tile_X0C_Y09_hi_out)
);
mantle_wire__typeBit8 Tile_X0C_Y09_lo (
    .in(Tile_X0C_Y09_lo_unq1),
    .out(Tile_X0C_Y09_lo_out)
);
wire [15:0] Tile_X0C_Y09_tile_id_out;
assign Tile_X0C_Y09_tile_id_out = {Tile_X0C_Y09_lo_out[7],Tile_X0C_Y09_lo_out[7:6],Tile_X0C_Y09_lo_out[6],Tile_X0C_Y09_hi_out[6:5],Tile_X0C_Y09_lo_out[4],Tile_X0C_Y09_lo_out[4:3],Tile_X0C_Y09_lo_out[3:2],Tile_X0C_Y09_lo_out[2],Tile_X0C_Y09_hi_out[2],Tile_X0C_Y09_lo_out[1:0],Tile_X0C_Y09_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X0C_Y09_tile_id (
    .in(Tile_X0C_Y09_tile_id_in),
    .out(Tile_X0C_Y09_tile_id_out)
);
Tile_PE Tile_X0C_Y0A (
    .SB_T0_EAST_SB_IN_B1(Tile_X0D_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0D_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0C_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0C_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0C_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0C_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0C_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0C_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0C_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0C_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0C_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0C_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0B_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0B_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0C_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0C_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0D_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0D_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0C_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0C_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0C_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0C_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0C_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0C_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0C_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0C_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0C_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0C_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0B_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0B_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0C_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0C_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0D_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0D_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0C_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0C_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0C_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0C_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0C_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0C_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0C_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0C_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0C_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0C_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0B_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0B_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0C_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0C_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0D_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0D_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0C_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0C_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0C_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0C_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0C_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0C_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0C_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0C_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0C_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0C_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0B_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0B_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0C_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0C_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0D_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0D_Y0A_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0C_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0C_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0C_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0C_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0C_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0C_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0C_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0C_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0C_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0C_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0B_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0B_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0C_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0C_Y0A_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0C_Y09_clk_out),
    .clk_out(Tile_X0C_Y0A_clk_out),
    .clk_pass_through(Tile_X0C_Y09_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0C_Y0A_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0C_Y0A_clk_pass_through_out_right),
    .config_config_addr(Tile_X0C_Y09_config_out_config_addr),
    .config_config_data(Tile_X0C_Y09_config_out_config_data),
    .config_out_config_addr(Tile_X0C_Y0A_config_out_config_addr),
    .config_out_config_data(Tile_X0C_Y0A_config_out_config_data),
    .config_out_read(Tile_X0C_Y0A_config_out_read),
    .config_out_write(Tile_X0C_Y0A_config_out_write),
    .config_read(Tile_X0C_Y09_config_out_read),
    .config_write(Tile_X0C_Y09_config_out_write),
    .hi(Tile_X0C_Y0A_hi_unq1),
    .lo(Tile_X0C_Y0A_lo_unq1),
    .read_config_data(Tile_X0C_Y0A_read_config_data),
    .read_config_data_in(Tile_X0C_Y09_read_config_data),
    .reset(Tile_X0C_Y09_reset_out),
    .reset_out(Tile_X0C_Y0A_reset_out),
    .stall(Tile_X0C_Y09_stall_out),
    .stall_out(Tile_X0C_Y0A_stall_out),
    .tile_id(Tile_X0C_Y0A_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0C_Y0A_hi (
    .in(Tile_X0C_Y0A_hi_unq1),
    .out(Tile_X0C_Y0A_hi_out)
);
mantle_wire__typeBit8 Tile_X0C_Y0A_lo (
    .in(Tile_X0C_Y0A_lo_unq1),
    .out(Tile_X0C_Y0A_lo_out)
);
wire [15:0] Tile_X0C_Y0A_tile_id_out;
assign Tile_X0C_Y0A_tile_id_out = {Tile_X0C_Y0A_lo_out[7],Tile_X0C_Y0A_lo_out[7:6],Tile_X0C_Y0A_lo_out[6],Tile_X0C_Y0A_hi_out[6:5],Tile_X0C_Y0A_lo_out[4],Tile_X0C_Y0A_lo_out[4:3],Tile_X0C_Y0A_lo_out[3:2],Tile_X0C_Y0A_lo_out[2],Tile_X0C_Y0A_hi_out[2],Tile_X0C_Y0A_lo_out[1],Tile_X0C_Y0A_hi_out[1],Tile_X0C_Y0A_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0C_Y0A_tile_id (
    .in(Tile_X0C_Y0A_tile_id_in),
    .out(Tile_X0C_Y0A_tile_id_out)
);
Tile_PE Tile_X0C_Y0B (
    .SB_T0_EAST_SB_IN_B1(Tile_X0D_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0D_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0C_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0C_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0C_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0C_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0C_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0C_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0C_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0C_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0C_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0C_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0B_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0B_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0C_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0C_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0D_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0D_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0C_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0C_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0C_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0C_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0C_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0C_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0C_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0C_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0C_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0C_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0B_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0B_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0C_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0C_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0D_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0D_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0C_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0C_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0C_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0C_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0C_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0C_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0C_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0C_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0C_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0C_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0B_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0B_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0C_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0C_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0D_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0D_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0C_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0C_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0C_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0C_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0C_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0C_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0C_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0C_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0C_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0C_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0B_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0B_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0C_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0C_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0D_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0D_Y0B_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0C_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0C_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0C_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0C_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0C_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0C_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0C_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0C_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0C_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0C_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0B_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0B_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0C_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0C_Y0B_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0C_Y0A_clk_out),
    .clk_out(Tile_X0C_Y0B_clk_out),
    .clk_pass_through(Tile_X0C_Y0A_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0C_Y0B_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0C_Y0B_clk_pass_through_out_right),
    .config_config_addr(Tile_X0C_Y0A_config_out_config_addr),
    .config_config_data(Tile_X0C_Y0A_config_out_config_data),
    .config_out_config_addr(Tile_X0C_Y0B_config_out_config_addr),
    .config_out_config_data(Tile_X0C_Y0B_config_out_config_data),
    .config_out_read(Tile_X0C_Y0B_config_out_read),
    .config_out_write(Tile_X0C_Y0B_config_out_write),
    .config_read(Tile_X0C_Y0A_config_out_read),
    .config_write(Tile_X0C_Y0A_config_out_write),
    .hi(Tile_X0C_Y0B_hi_unq1),
    .lo(Tile_X0C_Y0B_lo_unq1),
    .read_config_data(Tile_X0C_Y0B_read_config_data),
    .read_config_data_in(Tile_X0C_Y0A_read_config_data),
    .reset(Tile_X0C_Y0A_reset_out),
    .reset_out(Tile_X0C_Y0B_reset_out),
    .stall(Tile_X0C_Y0A_stall_out),
    .stall_out(Tile_X0C_Y0B_stall_out),
    .tile_id(Tile_X0C_Y0B_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0C_Y0B_hi (
    .in(Tile_X0C_Y0B_hi_unq1),
    .out(Tile_X0C_Y0B_hi_out)
);
mantle_wire__typeBit8 Tile_X0C_Y0B_lo (
    .in(Tile_X0C_Y0B_lo_unq1),
    .out(Tile_X0C_Y0B_lo_out)
);
wire [15:0] Tile_X0C_Y0B_tile_id_out;
assign Tile_X0C_Y0B_tile_id_out = {Tile_X0C_Y0B_lo_out[7],Tile_X0C_Y0B_lo_out[7:6],Tile_X0C_Y0B_lo_out[6],Tile_X0C_Y0B_hi_out[6:5],Tile_X0C_Y0B_lo_out[4],Tile_X0C_Y0B_lo_out[4:3],Tile_X0C_Y0B_lo_out[3:2],Tile_X0C_Y0B_lo_out[2],Tile_X0C_Y0B_hi_out[2],Tile_X0C_Y0B_lo_out[1],Tile_X0C_Y0B_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X0C_Y0B_tile_id (
    .in(Tile_X0C_Y0B_tile_id_in),
    .out(Tile_X0C_Y0B_tile_id_out)
);
Tile_PE Tile_X0C_Y0C (
    .SB_T0_EAST_SB_IN_B1(Tile_X0D_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0D_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0C_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0C_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0C_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0C_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0C_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0C_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0C_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0C_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0C_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0C_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0B_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0B_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0C_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0C_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0D_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0D_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0C_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0C_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0C_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0C_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0C_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0C_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0C_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0C_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0C_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0C_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0B_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0B_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0C_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0C_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0D_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0D_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0C_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0C_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0C_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0C_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0C_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0C_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0C_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0C_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0C_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0C_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0B_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0B_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0C_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0C_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0D_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0D_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0C_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0C_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0C_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0C_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0C_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0C_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0C_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0C_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0C_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0C_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0B_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0B_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0C_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0C_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0D_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0D_Y0C_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0C_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0C_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0C_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0C_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0C_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0C_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0C_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0C_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0C_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0C_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0B_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0B_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0C_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0C_Y0C_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0C_Y0B_clk_out),
    .clk_out(Tile_X0C_Y0C_clk_out),
    .clk_pass_through(Tile_X0C_Y0B_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0C_Y0C_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0C_Y0C_clk_pass_through_out_right),
    .config_config_addr(Tile_X0C_Y0B_config_out_config_addr),
    .config_config_data(Tile_X0C_Y0B_config_out_config_data),
    .config_out_config_addr(Tile_X0C_Y0C_config_out_config_addr),
    .config_out_config_data(Tile_X0C_Y0C_config_out_config_data),
    .config_out_read(Tile_X0C_Y0C_config_out_read),
    .config_out_write(Tile_X0C_Y0C_config_out_write),
    .config_read(Tile_X0C_Y0B_config_out_read),
    .config_write(Tile_X0C_Y0B_config_out_write),
    .hi(Tile_X0C_Y0C_hi_unq1),
    .lo(Tile_X0C_Y0C_lo_unq1),
    .read_config_data(Tile_X0C_Y0C_read_config_data),
    .read_config_data_in(Tile_X0C_Y0B_read_config_data),
    .reset(Tile_X0C_Y0B_reset_out),
    .reset_out(Tile_X0C_Y0C_reset_out),
    .stall(Tile_X0C_Y0B_stall_out),
    .stall_out(Tile_X0C_Y0C_stall_out),
    .tile_id(Tile_X0C_Y0C_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0C_Y0C_hi (
    .in(Tile_X0C_Y0C_hi_unq1),
    .out(Tile_X0C_Y0C_hi_out)
);
mantle_wire__typeBit8 Tile_X0C_Y0C_lo (
    .in(Tile_X0C_Y0C_lo_unq1),
    .out(Tile_X0C_Y0C_lo_out)
);
wire [15:0] Tile_X0C_Y0C_tile_id_out;
assign Tile_X0C_Y0C_tile_id_out = {Tile_X0C_Y0C_lo_out[7],Tile_X0C_Y0C_lo_out[7:6],Tile_X0C_Y0C_lo_out[6],Tile_X0C_Y0C_hi_out[6:5],Tile_X0C_Y0C_lo_out[4],Tile_X0C_Y0C_lo_out[4:3],Tile_X0C_Y0C_lo_out[3:2],Tile_X0C_Y0C_lo_out[2],Tile_X0C_Y0C_hi_out[2:1],Tile_X0C_Y0C_lo_out[0],Tile_X0C_Y0C_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0C_Y0C_tile_id (
    .in(Tile_X0C_Y0C_tile_id_in),
    .out(Tile_X0C_Y0C_tile_id_out)
);
Tile_PE Tile_X0C_Y0D (
    .SB_T0_EAST_SB_IN_B1(Tile_X0D_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0D_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0C_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0C_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0C_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0C_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0C_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0C_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0C_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0C_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0C_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0C_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0B_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0B_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0C_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0C_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0D_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0D_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0C_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0C_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0C_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0C_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0C_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0C_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0C_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0C_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0C_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0C_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0B_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0B_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0C_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0C_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0D_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0D_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0C_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0C_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0C_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0C_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0C_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0C_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0C_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0C_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0C_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0C_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0B_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0B_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0C_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0C_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0D_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0D_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0C_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0C_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0C_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0C_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0C_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0C_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0C_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0C_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0C_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0C_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0B_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0B_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0C_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0C_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0D_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0D_Y0D_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0C_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0C_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0C_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0C_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0C_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0C_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0C_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0C_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0C_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0C_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0B_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0B_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0C_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0C_Y0D_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0C_Y0C_clk_out),
    .clk_out(Tile_X0C_Y0D_clk_out),
    .clk_pass_through(Tile_X0C_Y0C_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0C_Y0D_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0C_Y0D_clk_pass_through_out_right),
    .config_config_addr(Tile_X0C_Y0C_config_out_config_addr),
    .config_config_data(Tile_X0C_Y0C_config_out_config_data),
    .config_out_config_addr(Tile_X0C_Y0D_config_out_config_addr),
    .config_out_config_data(Tile_X0C_Y0D_config_out_config_data),
    .config_out_read(Tile_X0C_Y0D_config_out_read),
    .config_out_write(Tile_X0C_Y0D_config_out_write),
    .config_read(Tile_X0C_Y0C_config_out_read),
    .config_write(Tile_X0C_Y0C_config_out_write),
    .hi(Tile_X0C_Y0D_hi_unq1),
    .lo(Tile_X0C_Y0D_lo_unq1),
    .read_config_data(Tile_X0C_Y0D_read_config_data),
    .read_config_data_in(Tile_X0C_Y0C_read_config_data),
    .reset(Tile_X0C_Y0C_reset_out),
    .reset_out(Tile_X0C_Y0D_reset_out),
    .stall(Tile_X0C_Y0C_stall_out),
    .stall_out(Tile_X0C_Y0D_stall_out),
    .tile_id(Tile_X0C_Y0D_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0C_Y0D_hi (
    .in(Tile_X0C_Y0D_hi_unq1),
    .out(Tile_X0C_Y0D_hi_out)
);
mantle_wire__typeBit8 Tile_X0C_Y0D_lo (
    .in(Tile_X0C_Y0D_lo_unq1),
    .out(Tile_X0C_Y0D_lo_out)
);
wire [15:0] Tile_X0C_Y0D_tile_id_out;
assign Tile_X0C_Y0D_tile_id_out = {Tile_X0C_Y0D_lo_out[7],Tile_X0C_Y0D_lo_out[7:6],Tile_X0C_Y0D_lo_out[6],Tile_X0C_Y0D_hi_out[6:5],Tile_X0C_Y0D_lo_out[4],Tile_X0C_Y0D_lo_out[4:3],Tile_X0C_Y0D_lo_out[3:2],Tile_X0C_Y0D_lo_out[2],Tile_X0C_Y0D_hi_out[2:1],Tile_X0C_Y0D_lo_out[0],Tile_X0C_Y0D_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X0C_Y0D_tile_id (
    .in(Tile_X0C_Y0D_tile_id_in),
    .out(Tile_X0C_Y0D_tile_id_out)
);
Tile_PE Tile_X0C_Y0E (
    .SB_T0_EAST_SB_IN_B1(Tile_X0D_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0D_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0C_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0C_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0C_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0C_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0C_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0C_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0C_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0C_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0C_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0C_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0B_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0B_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0C_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0C_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0D_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0D_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0C_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0C_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0C_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0C_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0C_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0C_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0C_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0C_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0C_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0C_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0B_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0B_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0C_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0C_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0D_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0D_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0C_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0C_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0C_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0C_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0C_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0C_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0C_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0C_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0C_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0C_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0B_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0B_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0C_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0C_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0D_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0D_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0C_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0C_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0C_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0C_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0C_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0C_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0C_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0C_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0C_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0C_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0B_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0B_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0C_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0C_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0D_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0D_Y0E_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0C_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0C_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0C_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0C_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0C_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0C_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0C_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0C_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0C_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0C_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0B_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0B_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0C_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0C_Y0E_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0C_Y0D_clk_out),
    .clk_out(Tile_X0C_Y0E_clk_out),
    .clk_pass_through(Tile_X0C_Y0D_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0C_Y0E_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0C_Y0E_clk_pass_through_out_right),
    .config_config_addr(Tile_X0C_Y0D_config_out_config_addr),
    .config_config_data(Tile_X0C_Y0D_config_out_config_data),
    .config_out_config_addr(Tile_X0C_Y0E_config_out_config_addr),
    .config_out_config_data(Tile_X0C_Y0E_config_out_config_data),
    .config_out_read(Tile_X0C_Y0E_config_out_read),
    .config_out_write(Tile_X0C_Y0E_config_out_write),
    .config_read(Tile_X0C_Y0D_config_out_read),
    .config_write(Tile_X0C_Y0D_config_out_write),
    .hi(Tile_X0C_Y0E_hi_unq1),
    .lo(Tile_X0C_Y0E_lo_unq1),
    .read_config_data(Tile_X0C_Y0E_read_config_data),
    .read_config_data_in(Tile_X0C_Y0D_read_config_data),
    .reset(Tile_X0C_Y0D_reset_out),
    .reset_out(Tile_X0C_Y0E_reset_out),
    .stall(Tile_X0C_Y0D_stall_out),
    .stall_out(Tile_X0C_Y0E_stall_out),
    .tile_id(Tile_X0C_Y0E_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0C_Y0E_hi (
    .in(Tile_X0C_Y0E_hi_unq1),
    .out(Tile_X0C_Y0E_hi_out)
);
mantle_wire__typeBit8 Tile_X0C_Y0E_lo (
    .in(Tile_X0C_Y0E_lo_unq1),
    .out(Tile_X0C_Y0E_lo_out)
);
wire [15:0] Tile_X0C_Y0E_tile_id_out;
assign Tile_X0C_Y0E_tile_id_out = {Tile_X0C_Y0E_lo_out[7],Tile_X0C_Y0E_lo_out[7:6],Tile_X0C_Y0E_lo_out[6],Tile_X0C_Y0E_hi_out[6:5],Tile_X0C_Y0E_lo_out[4],Tile_X0C_Y0E_lo_out[4:3],Tile_X0C_Y0E_lo_out[3:2],Tile_X0C_Y0E_lo_out[2],Tile_X0C_Y0E_hi_out[2:1],Tile_X0C_Y0E_hi_out[1],Tile_X0C_Y0E_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0C_Y0E_tile_id (
    .in(Tile_X0C_Y0E_tile_id_in),
    .out(Tile_X0C_Y0E_tile_id_out)
);
Tile_PE Tile_X0C_Y0F (
    .SB_T0_EAST_SB_IN_B1(Tile_X0D_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0D_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0C_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0C_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0C_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0C_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0C_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0C_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0C_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0C_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0C_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0C_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0B_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0B_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0C_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0C_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0D_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0D_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0C_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0C_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0C_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0C_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0C_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0C_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0C_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0C_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0C_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0C_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0B_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0B_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0C_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0C_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0D_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0D_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0C_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0C_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0C_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0C_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0C_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0C_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0C_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0C_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0C_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0C_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0B_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0B_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0C_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0C_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0D_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0D_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0C_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0C_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0C_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0C_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0C_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0C_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0C_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0C_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0C_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0C_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0B_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0B_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0C_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0C_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0D_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0D_Y0F_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0C_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0C_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0C_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0C_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0C_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0C_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0C_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0C_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0C_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0C_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0B_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0B_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0C_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0C_Y0F_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0C_Y0E_clk_out),
    .clk_out(Tile_X0C_Y0F_clk_out),
    .clk_pass_through(Tile_X0C_Y0E_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0C_Y0F_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0C_Y0F_clk_pass_through_out_right),
    .config_config_addr(Tile_X0C_Y0E_config_out_config_addr),
    .config_config_data(Tile_X0C_Y0E_config_out_config_data),
    .config_out_config_addr(Tile_X0C_Y0F_config_out_config_addr),
    .config_out_config_data(Tile_X0C_Y0F_config_out_config_data),
    .config_out_read(Tile_X0C_Y0F_config_out_read),
    .config_out_write(Tile_X0C_Y0F_config_out_write),
    .config_read(Tile_X0C_Y0E_config_out_read),
    .config_write(Tile_X0C_Y0E_config_out_write),
    .hi(Tile_X0C_Y0F_hi_unq1),
    .lo(Tile_X0C_Y0F_lo_unq1),
    .read_config_data(Tile_X0C_Y0F_read_config_data),
    .read_config_data_in(Tile_X0C_Y0E_read_config_data),
    .reset(Tile_X0C_Y0E_reset_out),
    .reset_out(Tile_X0C_Y0F_reset_out),
    .stall(Tile_X0C_Y0E_stall_out),
    .stall_out(Tile_X0C_Y0F_stall_out),
    .tile_id(Tile_X0C_Y0F_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0C_Y0F_hi (
    .in(Tile_X0C_Y0F_hi_unq1),
    .out(Tile_X0C_Y0F_hi_out)
);
mantle_wire__typeBit8 Tile_X0C_Y0F_lo (
    .in(Tile_X0C_Y0F_lo_unq1),
    .out(Tile_X0C_Y0F_lo_out)
);
wire [15:0] Tile_X0C_Y0F_tile_id_out;
assign Tile_X0C_Y0F_tile_id_out = {Tile_X0C_Y0F_lo_out[7],Tile_X0C_Y0F_lo_out[7:6],Tile_X0C_Y0F_lo_out[6],Tile_X0C_Y0F_hi_out[6:5],Tile_X0C_Y0F_lo_out[4],Tile_X0C_Y0F_lo_out[4:3],Tile_X0C_Y0F_lo_out[3:2],Tile_X0C_Y0F_lo_out[2],Tile_X0C_Y0F_hi_out[2:1],Tile_X0C_Y0F_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X0C_Y0F_tile_id (
    .in(Tile_X0C_Y0F_tile_id_in),
    .out(Tile_X0C_Y0F_tile_id_out)
);
Tile_PE Tile_X0C_Y10 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0D_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0D_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0C_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0C_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0C_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0C_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0C_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0C_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T0_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0C_Y10_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0C_Y10_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0B_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0B_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0C_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0C_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0D_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0D_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0C_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0C_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0C_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0C_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0C_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0C_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T1_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0C_Y10_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0C_Y10_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0B_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0B_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0C_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0C_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0D_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0D_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0C_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0C_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0C_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0C_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0C_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0C_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T2_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0C_Y10_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0C_Y10_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0B_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0B_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0C_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0C_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0D_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0D_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0C_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0C_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0C_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0C_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0C_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0C_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T3_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0C_Y10_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0C_Y10_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0B_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0B_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0C_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0C_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0D_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0D_Y10_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0C_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0C_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0C_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0C_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0C_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0C_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T4_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0C_Y10_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0C_Y10_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0B_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0B_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0C_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0C_Y10_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0C_Y0F_clk_out),
    .clk_out(Tile_X0C_Y10_clk_out),
    .clk_pass_through(Tile_X0C_Y0F_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0C_Y10_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0C_Y10_clk_pass_through_out_right),
    .config_config_addr(Tile_X0C_Y0F_config_out_config_addr),
    .config_config_data(Tile_X0C_Y0F_config_out_config_data),
    .config_out_config_addr(Tile_X0C_Y10_config_out_config_addr),
    .config_out_config_data(Tile_X0C_Y10_config_out_config_data),
    .config_out_read(Tile_X0C_Y10_config_out_read),
    .config_out_write(Tile_X0C_Y10_config_out_write),
    .config_read(Tile_X0C_Y0F_config_out_read),
    .config_write(Tile_X0C_Y0F_config_out_write),
    .hi(Tile_X0C_Y10_hi_unq1),
    .lo(Tile_X0C_Y10_lo_unq1),
    .read_config_data(Tile_X0C_Y10_read_config_data),
    .read_config_data_in(Tile_X0C_Y0F_read_config_data),
    .reset(Tile_X0C_Y0F_reset_out),
    .reset_out(Tile_X0C_Y10_reset_out),
    .stall(Tile_X0C_Y0F_stall_out),
    .stall_out(Tile_X0C_Y10_stall_out),
    .tile_id(Tile_X0C_Y10_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0C_Y10_hi (
    .in(Tile_X0C_Y10_hi_unq1),
    .out(Tile_X0C_Y10_hi_out)
);
mantle_wire__typeBit8 Tile_X0C_Y10_lo (
    .in(Tile_X0C_Y10_lo_unq1),
    .out(Tile_X0C_Y10_lo_out)
);
wire [15:0] Tile_X0C_Y10_tile_id_out;
assign Tile_X0C_Y10_tile_id_out = {Tile_X0C_Y10_lo_out[7],Tile_X0C_Y10_lo_out[7:6],Tile_X0C_Y10_lo_out[6],Tile_X0C_Y10_hi_out[6:5],Tile_X0C_Y10_lo_out[4],Tile_X0C_Y10_lo_out[4:3],Tile_X0C_Y10_lo_out[3:2],Tile_X0C_Y10_hi_out[2],Tile_X0C_Y10_lo_out[1],Tile_X0C_Y10_lo_out[1:0],Tile_X0C_Y10_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0C_Y10_tile_id (
    .in(Tile_X0C_Y10_tile_id_in),
    .out(Tile_X0C_Y10_tile_id_out)
);
wire [15:0] Tile_X0D_Y00_tile_id;
assign Tile_X0D_Y00_tile_id = {Tile_X0D_Y00_lo[7],Tile_X0D_Y00_lo[7:6],Tile_X0D_Y00_lo[6],Tile_X0D_Y00_hi[6:5],Tile_X0D_Y00_lo[4],Tile_X0D_Y00_hi[4],Tile_X0D_Y00_lo[3],Tile_X0D_Y00_lo[3:2],Tile_X0D_Y00_lo[2:1],Tile_X0D_Y00_lo[1:0],Tile_X0D_Y00_lo[0]};
Tile_io_core Tile_X0D_Y00 (
    .tile_id(Tile_X0D_Y00_tile_id),
    .glb2io_1(glb2io_1_X0D_Y00),
    .f2io_1(Tile_X0D_Y01_SB_T0_NORTH_SB_OUT_B1),
    .io2glb_1(Tile_X0D_Y00_io2glb_1),
    .io2f_1(Tile_X0D_Y00_io2f_1),
    .glb2io_16(glb2io_16_X0D_Y00),
    .f2io_16(Tile_X0D_Y01_SB_T0_NORTH_SB_OUT_B16),
    .io2glb_16(Tile_X0D_Y00_io2glb_16),
    .io2f_16(Tile_X0D_Y00_io2f_16),
    .hi(Tile_X0D_Y00_hi),
    .lo(Tile_X0D_Y00_lo)
);
Tile_PE Tile_X0D_Y01 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0E_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0E_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0D_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0D_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0D_Y00_io2f_1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0D_Y00_io2f_16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0D_Y01_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0D_Y01_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0D_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0D_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0D_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0D_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0C_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0C_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0D_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0D_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0E_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0E_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0D_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0D_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0D_Y00_io2f_1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0D_Y00_io2f_16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0D_Y01_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0D_Y01_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0D_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0D_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0D_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0D_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0C_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0C_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0D_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0D_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0E_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0E_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0D_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0D_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0D_Y00_io2f_1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0D_Y00_io2f_16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0D_Y01_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0D_Y01_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0D_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0D_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0D_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0D_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0C_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0C_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0D_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0D_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0E_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0E_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0D_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0D_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0D_Y00_io2f_1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0D_Y00_io2f_16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0D_Y01_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0D_Y01_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0D_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0D_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0D_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0D_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0C_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0C_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0D_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0D_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0E_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0E_Y01_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0D_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0D_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0D_Y00_io2f_1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0D_Y00_io2f_16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0D_Y01_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0D_Y01_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0D_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0D_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0D_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0D_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0C_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0C_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0D_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0D_Y01_SB_T4_WEST_SB_OUT_B16),
    .clk(clk),
    .clk_out(Tile_X0D_Y01_clk_out),
    .clk_pass_through(clk),
    .clk_pass_through_out_bot(Tile_X0D_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0D_Y01_clk_pass_through_out_right),
    .config_config_addr(config_13_config_addr),
    .config_config_data(config_13_config_data),
    .config_out_config_addr(Tile_X0D_Y01_config_out_config_addr),
    .config_out_config_data(Tile_X0D_Y01_config_out_config_data),
    .config_out_read(Tile_X0D_Y01_config_out_read),
    .config_out_write(Tile_X0D_Y01_config_out_write),
    .config_read(config_13_read),
    .config_write(config_13_write),
    .hi(Tile_X0D_Y01_hi_unq1),
    .lo(Tile_X0D_Y01_lo_unq1),
    .read_config_data(Tile_X0D_Y01_read_config_data),
    .read_config_data_in(const_0_32_out),
    .reset(reset),
    .reset_out(Tile_X0D_Y01_reset_out),
    .stall(stall[13]),
    .stall_out(Tile_X0D_Y01_stall_out),
    .tile_id(Tile_X0D_Y01_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0D_Y01_hi (
    .in(Tile_X0D_Y01_hi_unq1),
    .out(Tile_X0D_Y01_hi_out)
);
mantle_wire__typeBit8 Tile_X0D_Y01_lo (
    .in(Tile_X0D_Y01_lo_unq1),
    .out(Tile_X0D_Y01_lo_out)
);
wire [15:0] Tile_X0D_Y01_tile_id_out;
assign Tile_X0D_Y01_tile_id_out = {Tile_X0D_Y01_lo_out[7],Tile_X0D_Y01_lo_out[7:6],Tile_X0D_Y01_lo_out[6],Tile_X0D_Y01_hi_out[6:5],Tile_X0D_Y01_lo_out[4],Tile_X0D_Y01_hi_out[4],Tile_X0D_Y01_lo_out[3],Tile_X0D_Y01_lo_out[3:2],Tile_X0D_Y01_lo_out[2:1],Tile_X0D_Y01_lo_out[1:0],Tile_X0D_Y01_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X0D_Y01_tile_id (
    .in(Tile_X0D_Y01_tile_id_in),
    .out(Tile_X0D_Y01_tile_id_out)
);
Tile_PE Tile_X0D_Y02 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0E_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0E_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0D_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0D_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0D_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0D_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0D_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0D_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0D_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0D_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0D_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0D_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0C_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0C_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0D_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0D_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0E_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0E_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0D_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0D_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0D_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0D_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0D_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0D_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0D_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0D_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0D_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0D_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0C_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0C_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0D_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0D_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0E_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0E_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0D_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0D_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0D_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0D_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0D_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0D_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0D_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0D_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0D_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0D_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0C_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0C_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0D_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0D_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0E_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0E_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0D_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0D_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0D_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0D_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0D_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0D_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0D_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0D_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0D_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0D_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0C_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0C_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0D_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0D_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0E_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0E_Y02_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0D_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0D_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0D_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0D_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0D_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0D_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0D_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0D_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0D_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0D_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0C_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0C_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0D_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0D_Y02_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0D_Y01_clk_out),
    .clk_out(Tile_X0D_Y02_clk_out),
    .clk_pass_through(Tile_X0D_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0D_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0D_Y02_clk_pass_through_out_right),
    .config_config_addr(Tile_X0D_Y01_config_out_config_addr),
    .config_config_data(Tile_X0D_Y01_config_out_config_data),
    .config_out_config_addr(Tile_X0D_Y02_config_out_config_addr),
    .config_out_config_data(Tile_X0D_Y02_config_out_config_data),
    .config_out_read(Tile_X0D_Y02_config_out_read),
    .config_out_write(Tile_X0D_Y02_config_out_write),
    .config_read(Tile_X0D_Y01_config_out_read),
    .config_write(Tile_X0D_Y01_config_out_write),
    .hi(Tile_X0D_Y02_hi_unq1),
    .lo(Tile_X0D_Y02_lo_unq1),
    .read_config_data(Tile_X0D_Y02_read_config_data),
    .read_config_data_in(Tile_X0D_Y01_read_config_data),
    .reset(Tile_X0D_Y01_reset_out),
    .reset_out(Tile_X0D_Y02_reset_out),
    .stall(Tile_X0D_Y01_stall_out),
    .stall_out(Tile_X0D_Y02_stall_out),
    .tile_id(Tile_X0D_Y02_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0D_Y02_hi (
    .in(Tile_X0D_Y02_hi_unq1),
    .out(Tile_X0D_Y02_hi_out)
);
mantle_wire__typeBit8 Tile_X0D_Y02_lo (
    .in(Tile_X0D_Y02_lo_unq1),
    .out(Tile_X0D_Y02_lo_out)
);
wire [15:0] Tile_X0D_Y02_tile_id_out;
assign Tile_X0D_Y02_tile_id_out = {Tile_X0D_Y02_lo_out[7],Tile_X0D_Y02_lo_out[7:6],Tile_X0D_Y02_lo_out[6],Tile_X0D_Y02_hi_out[6:5],Tile_X0D_Y02_lo_out[4],Tile_X0D_Y02_hi_out[4],Tile_X0D_Y02_lo_out[3],Tile_X0D_Y02_lo_out[3:2],Tile_X0D_Y02_lo_out[2:1],Tile_X0D_Y02_lo_out[1],Tile_X0D_Y02_hi_out[1],Tile_X0D_Y02_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0D_Y02_tile_id (
    .in(Tile_X0D_Y02_tile_id_in),
    .out(Tile_X0D_Y02_tile_id_out)
);
Tile_PE Tile_X0D_Y03 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0E_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0E_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0D_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0D_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0D_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0D_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0D_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0D_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0D_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0D_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0D_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0D_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0C_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0C_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0D_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0D_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0E_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0E_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0D_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0D_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0D_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0D_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0D_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0D_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0D_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0D_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0D_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0D_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0C_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0C_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0D_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0D_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0E_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0E_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0D_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0D_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0D_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0D_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0D_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0D_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0D_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0D_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0D_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0D_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0C_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0C_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0D_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0D_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0E_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0E_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0D_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0D_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0D_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0D_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0D_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0D_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0D_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0D_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0D_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0D_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0C_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0C_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0D_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0D_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0E_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0E_Y03_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0D_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0D_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0D_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0D_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0D_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0D_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0D_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0D_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0D_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0D_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0C_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0C_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0D_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0D_Y03_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0D_Y02_clk_out),
    .clk_out(Tile_X0D_Y03_clk_out),
    .clk_pass_through(Tile_X0D_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0D_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0D_Y03_clk_pass_through_out_right),
    .config_config_addr(Tile_X0D_Y02_config_out_config_addr),
    .config_config_data(Tile_X0D_Y02_config_out_config_data),
    .config_out_config_addr(Tile_X0D_Y03_config_out_config_addr),
    .config_out_config_data(Tile_X0D_Y03_config_out_config_data),
    .config_out_read(Tile_X0D_Y03_config_out_read),
    .config_out_write(Tile_X0D_Y03_config_out_write),
    .config_read(Tile_X0D_Y02_config_out_read),
    .config_write(Tile_X0D_Y02_config_out_write),
    .hi(Tile_X0D_Y03_hi_unq1),
    .lo(Tile_X0D_Y03_lo_unq1),
    .read_config_data(Tile_X0D_Y03_read_config_data),
    .read_config_data_in(Tile_X0D_Y02_read_config_data),
    .reset(Tile_X0D_Y02_reset_out),
    .reset_out(Tile_X0D_Y03_reset_out),
    .stall(Tile_X0D_Y02_stall_out),
    .stall_out(Tile_X0D_Y03_stall_out),
    .tile_id(Tile_X0D_Y03_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0D_Y03_hi (
    .in(Tile_X0D_Y03_hi_unq1),
    .out(Tile_X0D_Y03_hi_out)
);
mantle_wire__typeBit8 Tile_X0D_Y03_lo (
    .in(Tile_X0D_Y03_lo_unq1),
    .out(Tile_X0D_Y03_lo_out)
);
wire [15:0] Tile_X0D_Y03_tile_id_out;
assign Tile_X0D_Y03_tile_id_out = {Tile_X0D_Y03_lo_out[7],Tile_X0D_Y03_lo_out[7:6],Tile_X0D_Y03_lo_out[6],Tile_X0D_Y03_hi_out[6:5],Tile_X0D_Y03_lo_out[4],Tile_X0D_Y03_hi_out[4],Tile_X0D_Y03_lo_out[3],Tile_X0D_Y03_lo_out[3:2],Tile_X0D_Y03_lo_out[2:1],Tile_X0D_Y03_lo_out[1],Tile_X0D_Y03_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X0D_Y03_tile_id (
    .in(Tile_X0D_Y03_tile_id_in),
    .out(Tile_X0D_Y03_tile_id_out)
);
Tile_PE Tile_X0D_Y04 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0E_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0E_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0D_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0D_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0D_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0D_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0D_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0D_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0D_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0D_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0D_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0D_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0C_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0C_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0D_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0D_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0E_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0E_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0D_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0D_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0D_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0D_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0D_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0D_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0D_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0D_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0D_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0D_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0C_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0C_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0D_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0D_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0E_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0E_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0D_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0D_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0D_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0D_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0D_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0D_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0D_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0D_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0D_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0D_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0C_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0C_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0D_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0D_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0E_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0E_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0D_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0D_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0D_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0D_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0D_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0D_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0D_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0D_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0D_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0D_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0C_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0C_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0D_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0D_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0E_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0E_Y04_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0D_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0D_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0D_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0D_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0D_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0D_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0D_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0D_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0D_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0D_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0C_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0C_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0D_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0D_Y04_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0D_Y03_clk_out),
    .clk_out(Tile_X0D_Y04_clk_out),
    .clk_pass_through(Tile_X0D_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0D_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0D_Y04_clk_pass_through_out_right),
    .config_config_addr(Tile_X0D_Y03_config_out_config_addr),
    .config_config_data(Tile_X0D_Y03_config_out_config_data),
    .config_out_config_addr(Tile_X0D_Y04_config_out_config_addr),
    .config_out_config_data(Tile_X0D_Y04_config_out_config_data),
    .config_out_read(Tile_X0D_Y04_config_out_read),
    .config_out_write(Tile_X0D_Y04_config_out_write),
    .config_read(Tile_X0D_Y03_config_out_read),
    .config_write(Tile_X0D_Y03_config_out_write),
    .hi(Tile_X0D_Y04_hi_unq1),
    .lo(Tile_X0D_Y04_lo_unq1),
    .read_config_data(Tile_X0D_Y04_read_config_data),
    .read_config_data_in(Tile_X0D_Y03_read_config_data),
    .reset(Tile_X0D_Y03_reset_out),
    .reset_out(Tile_X0D_Y04_reset_out),
    .stall(Tile_X0D_Y03_stall_out),
    .stall_out(Tile_X0D_Y04_stall_out),
    .tile_id(Tile_X0D_Y04_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0D_Y04_hi (
    .in(Tile_X0D_Y04_hi_unq1),
    .out(Tile_X0D_Y04_hi_out)
);
mantle_wire__typeBit8 Tile_X0D_Y04_lo (
    .in(Tile_X0D_Y04_lo_unq1),
    .out(Tile_X0D_Y04_lo_out)
);
wire [15:0] Tile_X0D_Y04_tile_id_out;
assign Tile_X0D_Y04_tile_id_out = {Tile_X0D_Y04_lo_out[7],Tile_X0D_Y04_lo_out[7:6],Tile_X0D_Y04_lo_out[6],Tile_X0D_Y04_hi_out[6:5],Tile_X0D_Y04_lo_out[4],Tile_X0D_Y04_hi_out[4],Tile_X0D_Y04_lo_out[3],Tile_X0D_Y04_lo_out[3:2],Tile_X0D_Y04_lo_out[2:1],Tile_X0D_Y04_hi_out[1],Tile_X0D_Y04_lo_out[0],Tile_X0D_Y04_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0D_Y04_tile_id (
    .in(Tile_X0D_Y04_tile_id_in),
    .out(Tile_X0D_Y04_tile_id_out)
);
Tile_PE Tile_X0D_Y05 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0E_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0E_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0D_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0D_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0D_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0D_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0D_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0D_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0D_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0D_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0D_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0D_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0C_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0C_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0D_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0D_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0E_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0E_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0D_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0D_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0D_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0D_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0D_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0D_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0D_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0D_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0D_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0D_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0C_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0C_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0D_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0D_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0E_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0E_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0D_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0D_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0D_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0D_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0D_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0D_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0D_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0D_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0D_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0D_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0C_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0C_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0D_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0D_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0E_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0E_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0D_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0D_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0D_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0D_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0D_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0D_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0D_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0D_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0D_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0D_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0C_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0C_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0D_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0D_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0E_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0E_Y05_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0D_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0D_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0D_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0D_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0D_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0D_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0D_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0D_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0D_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0D_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0C_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0C_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0D_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0D_Y05_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0D_Y04_clk_out),
    .clk_out(Tile_X0D_Y05_clk_out),
    .clk_pass_through(Tile_X0D_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0D_Y05_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0D_Y05_clk_pass_through_out_right),
    .config_config_addr(Tile_X0D_Y04_config_out_config_addr),
    .config_config_data(Tile_X0D_Y04_config_out_config_data),
    .config_out_config_addr(Tile_X0D_Y05_config_out_config_addr),
    .config_out_config_data(Tile_X0D_Y05_config_out_config_data),
    .config_out_read(Tile_X0D_Y05_config_out_read),
    .config_out_write(Tile_X0D_Y05_config_out_write),
    .config_read(Tile_X0D_Y04_config_out_read),
    .config_write(Tile_X0D_Y04_config_out_write),
    .hi(Tile_X0D_Y05_hi_unq1),
    .lo(Tile_X0D_Y05_lo_unq1),
    .read_config_data(Tile_X0D_Y05_read_config_data),
    .read_config_data_in(Tile_X0D_Y04_read_config_data),
    .reset(Tile_X0D_Y04_reset_out),
    .reset_out(Tile_X0D_Y05_reset_out),
    .stall(Tile_X0D_Y04_stall_out),
    .stall_out(Tile_X0D_Y05_stall_out),
    .tile_id(Tile_X0D_Y05_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0D_Y05_hi (
    .in(Tile_X0D_Y05_hi_unq1),
    .out(Tile_X0D_Y05_hi_out)
);
mantle_wire__typeBit8 Tile_X0D_Y05_lo (
    .in(Tile_X0D_Y05_lo_unq1),
    .out(Tile_X0D_Y05_lo_out)
);
wire [15:0] Tile_X0D_Y05_tile_id_out;
assign Tile_X0D_Y05_tile_id_out = {Tile_X0D_Y05_lo_out[7],Tile_X0D_Y05_lo_out[7:6],Tile_X0D_Y05_lo_out[6],Tile_X0D_Y05_hi_out[6:5],Tile_X0D_Y05_lo_out[4],Tile_X0D_Y05_hi_out[4],Tile_X0D_Y05_lo_out[3],Tile_X0D_Y05_lo_out[3:2],Tile_X0D_Y05_lo_out[2:1],Tile_X0D_Y05_hi_out[1],Tile_X0D_Y05_lo_out[0],Tile_X0D_Y05_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X0D_Y05_tile_id (
    .in(Tile_X0D_Y05_tile_id_in),
    .out(Tile_X0D_Y05_tile_id_out)
);
Tile_PE Tile_X0D_Y06 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0E_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0E_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0D_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0D_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0D_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0D_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0D_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0D_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0D_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0D_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0D_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0D_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0C_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0C_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0D_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0D_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0E_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0E_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0D_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0D_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0D_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0D_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0D_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0D_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0D_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0D_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0D_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0D_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0C_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0C_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0D_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0D_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0E_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0E_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0D_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0D_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0D_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0D_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0D_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0D_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0D_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0D_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0D_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0D_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0C_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0C_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0D_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0D_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0E_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0E_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0D_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0D_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0D_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0D_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0D_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0D_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0D_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0D_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0D_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0D_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0C_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0C_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0D_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0D_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0E_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0E_Y06_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0D_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0D_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0D_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0D_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0D_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0D_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0D_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0D_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0D_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0D_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0C_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0C_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0D_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0D_Y06_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0D_Y05_clk_out),
    .clk_out(Tile_X0D_Y06_clk_out),
    .clk_pass_through(Tile_X0D_Y05_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0D_Y06_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0D_Y06_clk_pass_through_out_right),
    .config_config_addr(Tile_X0D_Y05_config_out_config_addr),
    .config_config_data(Tile_X0D_Y05_config_out_config_data),
    .config_out_config_addr(Tile_X0D_Y06_config_out_config_addr),
    .config_out_config_data(Tile_X0D_Y06_config_out_config_data),
    .config_out_read(Tile_X0D_Y06_config_out_read),
    .config_out_write(Tile_X0D_Y06_config_out_write),
    .config_read(Tile_X0D_Y05_config_out_read),
    .config_write(Tile_X0D_Y05_config_out_write),
    .hi(Tile_X0D_Y06_hi_unq1),
    .lo(Tile_X0D_Y06_lo_unq1),
    .read_config_data(Tile_X0D_Y06_read_config_data),
    .read_config_data_in(Tile_X0D_Y05_read_config_data),
    .reset(Tile_X0D_Y05_reset_out),
    .reset_out(Tile_X0D_Y06_reset_out),
    .stall(Tile_X0D_Y05_stall_out),
    .stall_out(Tile_X0D_Y06_stall_out),
    .tile_id(Tile_X0D_Y06_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0D_Y06_hi (
    .in(Tile_X0D_Y06_hi_unq1),
    .out(Tile_X0D_Y06_hi_out)
);
mantle_wire__typeBit8 Tile_X0D_Y06_lo (
    .in(Tile_X0D_Y06_lo_unq1),
    .out(Tile_X0D_Y06_lo_out)
);
wire [15:0] Tile_X0D_Y06_tile_id_out;
assign Tile_X0D_Y06_tile_id_out = {Tile_X0D_Y06_lo_out[7],Tile_X0D_Y06_lo_out[7:6],Tile_X0D_Y06_lo_out[6],Tile_X0D_Y06_hi_out[6:5],Tile_X0D_Y06_lo_out[4],Tile_X0D_Y06_hi_out[4],Tile_X0D_Y06_lo_out[3],Tile_X0D_Y06_lo_out[3:2],Tile_X0D_Y06_lo_out[2:1],Tile_X0D_Y06_hi_out[1],Tile_X0D_Y06_hi_out[1],Tile_X0D_Y06_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0D_Y06_tile_id (
    .in(Tile_X0D_Y06_tile_id_in),
    .out(Tile_X0D_Y06_tile_id_out)
);
Tile_PE Tile_X0D_Y07 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0E_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0E_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0D_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0D_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0D_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0D_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0D_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0D_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0D_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0D_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0D_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0D_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0C_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0C_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0D_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0D_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0E_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0E_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0D_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0D_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0D_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0D_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0D_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0D_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0D_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0D_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0D_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0D_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0C_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0C_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0D_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0D_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0E_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0E_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0D_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0D_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0D_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0D_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0D_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0D_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0D_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0D_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0D_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0D_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0C_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0C_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0D_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0D_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0E_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0E_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0D_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0D_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0D_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0D_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0D_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0D_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0D_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0D_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0D_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0D_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0C_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0C_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0D_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0D_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0E_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0E_Y07_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0D_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0D_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0D_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0D_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0D_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0D_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0D_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0D_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0D_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0D_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0C_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0C_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0D_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0D_Y07_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0D_Y06_clk_out),
    .clk_out(Tile_X0D_Y07_clk_out),
    .clk_pass_through(Tile_X0D_Y06_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0D_Y07_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0D_Y07_clk_pass_through_out_right),
    .config_config_addr(Tile_X0D_Y06_config_out_config_addr),
    .config_config_data(Tile_X0D_Y06_config_out_config_data),
    .config_out_config_addr(Tile_X0D_Y07_config_out_config_addr),
    .config_out_config_data(Tile_X0D_Y07_config_out_config_data),
    .config_out_read(Tile_X0D_Y07_config_out_read),
    .config_out_write(Tile_X0D_Y07_config_out_write),
    .config_read(Tile_X0D_Y06_config_out_read),
    .config_write(Tile_X0D_Y06_config_out_write),
    .hi(Tile_X0D_Y07_hi_unq1),
    .lo(Tile_X0D_Y07_lo_unq1),
    .read_config_data(Tile_X0D_Y07_read_config_data),
    .read_config_data_in(Tile_X0D_Y06_read_config_data),
    .reset(Tile_X0D_Y06_reset_out),
    .reset_out(Tile_X0D_Y07_reset_out),
    .stall(Tile_X0D_Y06_stall_out),
    .stall_out(Tile_X0D_Y07_stall_out),
    .tile_id(Tile_X0D_Y07_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0D_Y07_hi (
    .in(Tile_X0D_Y07_hi_unq1),
    .out(Tile_X0D_Y07_hi_out)
);
mantle_wire__typeBit8 Tile_X0D_Y07_lo (
    .in(Tile_X0D_Y07_lo_unq1),
    .out(Tile_X0D_Y07_lo_out)
);
wire [15:0] Tile_X0D_Y07_tile_id_out;
assign Tile_X0D_Y07_tile_id_out = {Tile_X0D_Y07_lo_out[7],Tile_X0D_Y07_lo_out[7:6],Tile_X0D_Y07_lo_out[6],Tile_X0D_Y07_hi_out[6:5],Tile_X0D_Y07_lo_out[4],Tile_X0D_Y07_hi_out[4],Tile_X0D_Y07_lo_out[3],Tile_X0D_Y07_lo_out[3:2],Tile_X0D_Y07_lo_out[2:1],Tile_X0D_Y07_hi_out[1],Tile_X0D_Y07_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X0D_Y07_tile_id (
    .in(Tile_X0D_Y07_tile_id_in),
    .out(Tile_X0D_Y07_tile_id_out)
);
Tile_PE Tile_X0D_Y08 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0E_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0E_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0D_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0D_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0D_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0D_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0D_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0D_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0D_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0D_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0D_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0D_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0C_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0C_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0D_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0D_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0E_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0E_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0D_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0D_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0D_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0D_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0D_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0D_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0D_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0D_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0D_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0D_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0C_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0C_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0D_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0D_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0E_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0E_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0D_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0D_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0D_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0D_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0D_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0D_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0D_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0D_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0D_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0D_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0C_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0C_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0D_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0D_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0E_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0E_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0D_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0D_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0D_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0D_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0D_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0D_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0D_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0D_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0D_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0D_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0C_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0C_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0D_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0D_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0E_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0E_Y08_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0D_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0D_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0D_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0D_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0D_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0D_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0D_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0D_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0D_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0D_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0C_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0C_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0D_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0D_Y08_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0D_Y07_clk_out),
    .clk_out(Tile_X0D_Y08_clk_out),
    .clk_pass_through(Tile_X0D_Y07_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0D_Y08_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0D_Y08_clk_pass_through_out_right),
    .config_config_addr(Tile_X0D_Y07_config_out_config_addr),
    .config_config_data(Tile_X0D_Y07_config_out_config_data),
    .config_out_config_addr(Tile_X0D_Y08_config_out_config_addr),
    .config_out_config_data(Tile_X0D_Y08_config_out_config_data),
    .config_out_read(Tile_X0D_Y08_config_out_read),
    .config_out_write(Tile_X0D_Y08_config_out_write),
    .config_read(Tile_X0D_Y07_config_out_read),
    .config_write(Tile_X0D_Y07_config_out_write),
    .hi(Tile_X0D_Y08_hi_unq1),
    .lo(Tile_X0D_Y08_lo_unq1),
    .read_config_data(Tile_X0D_Y08_read_config_data),
    .read_config_data_in(Tile_X0D_Y07_read_config_data),
    .reset(Tile_X0D_Y07_reset_out),
    .reset_out(Tile_X0D_Y08_reset_out),
    .stall(Tile_X0D_Y07_stall_out),
    .stall_out(Tile_X0D_Y08_stall_out),
    .tile_id(Tile_X0D_Y08_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0D_Y08_hi (
    .in(Tile_X0D_Y08_hi_unq1),
    .out(Tile_X0D_Y08_hi_out)
);
mantle_wire__typeBit8 Tile_X0D_Y08_lo (
    .in(Tile_X0D_Y08_lo_unq1),
    .out(Tile_X0D_Y08_lo_out)
);
wire [15:0] Tile_X0D_Y08_tile_id_out;
assign Tile_X0D_Y08_tile_id_out = {Tile_X0D_Y08_lo_out[7],Tile_X0D_Y08_lo_out[7:6],Tile_X0D_Y08_lo_out[6],Tile_X0D_Y08_hi_out[6:5],Tile_X0D_Y08_lo_out[4],Tile_X0D_Y08_hi_out[4],Tile_X0D_Y08_lo_out[3],Tile_X0D_Y08_lo_out[3:2],Tile_X0D_Y08_lo_out[2],Tile_X0D_Y08_hi_out[2],Tile_X0D_Y08_lo_out[1:0],Tile_X0D_Y08_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0D_Y08_tile_id (
    .in(Tile_X0D_Y08_tile_id_in),
    .out(Tile_X0D_Y08_tile_id_out)
);
Tile_PE Tile_X0D_Y09 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0E_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0E_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0D_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0D_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0D_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0D_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0D_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0D_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0D_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0D_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0D_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0D_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0C_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0C_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0D_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0D_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0E_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0E_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0D_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0D_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0D_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0D_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0D_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0D_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0D_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0D_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0D_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0D_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0C_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0C_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0D_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0D_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0E_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0E_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0D_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0D_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0D_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0D_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0D_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0D_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0D_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0D_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0D_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0D_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0C_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0C_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0D_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0D_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0E_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0E_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0D_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0D_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0D_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0D_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0D_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0D_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0D_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0D_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0D_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0D_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0C_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0C_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0D_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0D_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0E_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0E_Y09_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0D_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0D_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0D_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0D_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0D_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0D_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0D_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0D_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0D_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0D_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0C_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0C_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0D_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0D_Y09_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0D_Y08_clk_out),
    .clk_out(Tile_X0D_Y09_clk_out),
    .clk_pass_through(Tile_X0D_Y08_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0D_Y09_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0D_Y09_clk_pass_through_out_right),
    .config_config_addr(ConfigPipeStage_inst13_config_out_config_addr),
    .config_config_data(ConfigPipeStage_inst13_config_out_config_data),
    .config_out_config_addr(Tile_X0D_Y09_config_out_config_addr),
    .config_out_config_data(Tile_X0D_Y09_config_out_config_data),
    .config_out_read(Tile_X0D_Y09_config_out_read),
    .config_out_write(Tile_X0D_Y09_config_out_write),
    .config_read(ConfigPipeStage_inst13_config_out_read),
    .config_write(ConfigPipeStage_inst13_config_out_write),
    .hi(Tile_X0D_Y09_hi_unq1),
    .lo(Tile_X0D_Y09_lo_unq1),
    .read_config_data(Tile_X0D_Y09_read_config_data),
    .read_config_data_in(Tile_X0D_Y08_read_config_data),
    .reset(Tile_X0D_Y08_reset_out),
    .reset_out(Tile_X0D_Y09_reset_out),
    .stall(Tile_X0D_Y08_stall_out),
    .stall_out(Tile_X0D_Y09_stall_out),
    .tile_id(Tile_X0D_Y09_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0D_Y09_hi (
    .in(Tile_X0D_Y09_hi_unq1),
    .out(Tile_X0D_Y09_hi_out)
);
mantle_wire__typeBit8 Tile_X0D_Y09_lo (
    .in(Tile_X0D_Y09_lo_unq1),
    .out(Tile_X0D_Y09_lo_out)
);
wire [15:0] Tile_X0D_Y09_tile_id_out;
assign Tile_X0D_Y09_tile_id_out = {Tile_X0D_Y09_lo_out[7],Tile_X0D_Y09_lo_out[7:6],Tile_X0D_Y09_lo_out[6],Tile_X0D_Y09_hi_out[6:5],Tile_X0D_Y09_lo_out[4],Tile_X0D_Y09_hi_out[4],Tile_X0D_Y09_lo_out[3],Tile_X0D_Y09_lo_out[3:2],Tile_X0D_Y09_lo_out[2],Tile_X0D_Y09_hi_out[2],Tile_X0D_Y09_lo_out[1:0],Tile_X0D_Y09_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X0D_Y09_tile_id (
    .in(Tile_X0D_Y09_tile_id_in),
    .out(Tile_X0D_Y09_tile_id_out)
);
Tile_PE Tile_X0D_Y0A (
    .SB_T0_EAST_SB_IN_B1(Tile_X0E_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0E_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0D_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0D_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0D_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0D_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0D_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0D_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0D_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0D_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0D_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0D_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0C_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0C_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0D_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0D_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0E_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0E_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0D_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0D_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0D_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0D_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0D_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0D_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0D_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0D_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0D_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0D_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0C_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0C_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0D_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0D_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0E_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0E_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0D_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0D_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0D_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0D_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0D_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0D_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0D_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0D_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0D_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0D_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0C_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0C_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0D_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0D_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0E_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0E_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0D_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0D_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0D_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0D_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0D_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0D_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0D_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0D_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0D_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0D_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0C_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0C_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0D_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0D_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0E_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0E_Y0A_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0D_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0D_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0D_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0D_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0D_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0D_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0D_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0D_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0D_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0D_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0C_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0C_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0D_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0D_Y0A_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0D_Y09_clk_out),
    .clk_out(Tile_X0D_Y0A_clk_out),
    .clk_pass_through(Tile_X0D_Y09_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0D_Y0A_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0D_Y0A_clk_pass_through_out_right),
    .config_config_addr(Tile_X0D_Y09_config_out_config_addr),
    .config_config_data(Tile_X0D_Y09_config_out_config_data),
    .config_out_config_addr(Tile_X0D_Y0A_config_out_config_addr),
    .config_out_config_data(Tile_X0D_Y0A_config_out_config_data),
    .config_out_read(Tile_X0D_Y0A_config_out_read),
    .config_out_write(Tile_X0D_Y0A_config_out_write),
    .config_read(Tile_X0D_Y09_config_out_read),
    .config_write(Tile_X0D_Y09_config_out_write),
    .hi(Tile_X0D_Y0A_hi_unq1),
    .lo(Tile_X0D_Y0A_lo_unq1),
    .read_config_data(Tile_X0D_Y0A_read_config_data),
    .read_config_data_in(Tile_X0D_Y09_read_config_data),
    .reset(Tile_X0D_Y09_reset_out),
    .reset_out(Tile_X0D_Y0A_reset_out),
    .stall(Tile_X0D_Y09_stall_out),
    .stall_out(Tile_X0D_Y0A_stall_out),
    .tile_id(Tile_X0D_Y0A_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0D_Y0A_hi (
    .in(Tile_X0D_Y0A_hi_unq1),
    .out(Tile_X0D_Y0A_hi_out)
);
mantle_wire__typeBit8 Tile_X0D_Y0A_lo (
    .in(Tile_X0D_Y0A_lo_unq1),
    .out(Tile_X0D_Y0A_lo_out)
);
wire [15:0] Tile_X0D_Y0A_tile_id_out;
assign Tile_X0D_Y0A_tile_id_out = {Tile_X0D_Y0A_lo_out[7],Tile_X0D_Y0A_lo_out[7:6],Tile_X0D_Y0A_lo_out[6],Tile_X0D_Y0A_hi_out[6:5],Tile_X0D_Y0A_lo_out[4],Tile_X0D_Y0A_hi_out[4],Tile_X0D_Y0A_lo_out[3],Tile_X0D_Y0A_lo_out[3:2],Tile_X0D_Y0A_lo_out[2],Tile_X0D_Y0A_hi_out[2],Tile_X0D_Y0A_lo_out[1],Tile_X0D_Y0A_hi_out[1],Tile_X0D_Y0A_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0D_Y0A_tile_id (
    .in(Tile_X0D_Y0A_tile_id_in),
    .out(Tile_X0D_Y0A_tile_id_out)
);
Tile_PE Tile_X0D_Y0B (
    .SB_T0_EAST_SB_IN_B1(Tile_X0E_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0E_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0D_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0D_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0D_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0D_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0D_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0D_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0D_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0D_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0D_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0D_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0C_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0C_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0D_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0D_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0E_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0E_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0D_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0D_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0D_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0D_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0D_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0D_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0D_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0D_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0D_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0D_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0C_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0C_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0D_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0D_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0E_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0E_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0D_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0D_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0D_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0D_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0D_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0D_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0D_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0D_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0D_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0D_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0C_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0C_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0D_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0D_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0E_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0E_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0D_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0D_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0D_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0D_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0D_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0D_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0D_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0D_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0D_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0D_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0C_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0C_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0D_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0D_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0E_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0E_Y0B_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0D_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0D_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0D_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0D_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0D_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0D_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0D_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0D_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0D_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0D_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0C_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0C_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0D_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0D_Y0B_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0D_Y0A_clk_out),
    .clk_out(Tile_X0D_Y0B_clk_out),
    .clk_pass_through(Tile_X0D_Y0A_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0D_Y0B_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0D_Y0B_clk_pass_through_out_right),
    .config_config_addr(Tile_X0D_Y0A_config_out_config_addr),
    .config_config_data(Tile_X0D_Y0A_config_out_config_data),
    .config_out_config_addr(Tile_X0D_Y0B_config_out_config_addr),
    .config_out_config_data(Tile_X0D_Y0B_config_out_config_data),
    .config_out_read(Tile_X0D_Y0B_config_out_read),
    .config_out_write(Tile_X0D_Y0B_config_out_write),
    .config_read(Tile_X0D_Y0A_config_out_read),
    .config_write(Tile_X0D_Y0A_config_out_write),
    .hi(Tile_X0D_Y0B_hi_unq1),
    .lo(Tile_X0D_Y0B_lo_unq1),
    .read_config_data(Tile_X0D_Y0B_read_config_data),
    .read_config_data_in(Tile_X0D_Y0A_read_config_data),
    .reset(Tile_X0D_Y0A_reset_out),
    .reset_out(Tile_X0D_Y0B_reset_out),
    .stall(Tile_X0D_Y0A_stall_out),
    .stall_out(Tile_X0D_Y0B_stall_out),
    .tile_id(Tile_X0D_Y0B_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0D_Y0B_hi (
    .in(Tile_X0D_Y0B_hi_unq1),
    .out(Tile_X0D_Y0B_hi_out)
);
mantle_wire__typeBit8 Tile_X0D_Y0B_lo (
    .in(Tile_X0D_Y0B_lo_unq1),
    .out(Tile_X0D_Y0B_lo_out)
);
wire [15:0] Tile_X0D_Y0B_tile_id_out;
assign Tile_X0D_Y0B_tile_id_out = {Tile_X0D_Y0B_lo_out[7],Tile_X0D_Y0B_lo_out[7:6],Tile_X0D_Y0B_lo_out[6],Tile_X0D_Y0B_hi_out[6:5],Tile_X0D_Y0B_lo_out[4],Tile_X0D_Y0B_hi_out[4],Tile_X0D_Y0B_lo_out[3],Tile_X0D_Y0B_lo_out[3:2],Tile_X0D_Y0B_lo_out[2],Tile_X0D_Y0B_hi_out[2],Tile_X0D_Y0B_lo_out[1],Tile_X0D_Y0B_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X0D_Y0B_tile_id (
    .in(Tile_X0D_Y0B_tile_id_in),
    .out(Tile_X0D_Y0B_tile_id_out)
);
Tile_PE Tile_X0D_Y0C (
    .SB_T0_EAST_SB_IN_B1(Tile_X0E_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0E_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0D_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0D_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0D_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0D_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0D_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0D_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0D_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0D_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0D_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0D_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0C_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0C_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0D_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0D_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0E_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0E_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0D_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0D_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0D_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0D_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0D_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0D_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0D_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0D_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0D_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0D_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0C_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0C_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0D_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0D_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0E_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0E_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0D_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0D_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0D_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0D_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0D_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0D_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0D_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0D_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0D_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0D_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0C_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0C_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0D_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0D_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0E_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0E_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0D_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0D_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0D_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0D_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0D_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0D_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0D_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0D_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0D_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0D_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0C_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0C_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0D_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0D_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0E_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0E_Y0C_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0D_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0D_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0D_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0D_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0D_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0D_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0D_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0D_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0D_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0D_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0C_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0C_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0D_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0D_Y0C_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0D_Y0B_clk_out),
    .clk_out(Tile_X0D_Y0C_clk_out),
    .clk_pass_through(Tile_X0D_Y0B_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0D_Y0C_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0D_Y0C_clk_pass_through_out_right),
    .config_config_addr(Tile_X0D_Y0B_config_out_config_addr),
    .config_config_data(Tile_X0D_Y0B_config_out_config_data),
    .config_out_config_addr(Tile_X0D_Y0C_config_out_config_addr),
    .config_out_config_data(Tile_X0D_Y0C_config_out_config_data),
    .config_out_read(Tile_X0D_Y0C_config_out_read),
    .config_out_write(Tile_X0D_Y0C_config_out_write),
    .config_read(Tile_X0D_Y0B_config_out_read),
    .config_write(Tile_X0D_Y0B_config_out_write),
    .hi(Tile_X0D_Y0C_hi_unq1),
    .lo(Tile_X0D_Y0C_lo_unq1),
    .read_config_data(Tile_X0D_Y0C_read_config_data),
    .read_config_data_in(Tile_X0D_Y0B_read_config_data),
    .reset(Tile_X0D_Y0B_reset_out),
    .reset_out(Tile_X0D_Y0C_reset_out),
    .stall(Tile_X0D_Y0B_stall_out),
    .stall_out(Tile_X0D_Y0C_stall_out),
    .tile_id(Tile_X0D_Y0C_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0D_Y0C_hi (
    .in(Tile_X0D_Y0C_hi_unq1),
    .out(Tile_X0D_Y0C_hi_out)
);
mantle_wire__typeBit8 Tile_X0D_Y0C_lo (
    .in(Tile_X0D_Y0C_lo_unq1),
    .out(Tile_X0D_Y0C_lo_out)
);
wire [15:0] Tile_X0D_Y0C_tile_id_out;
assign Tile_X0D_Y0C_tile_id_out = {Tile_X0D_Y0C_lo_out[7],Tile_X0D_Y0C_lo_out[7:6],Tile_X0D_Y0C_lo_out[6],Tile_X0D_Y0C_hi_out[6:5],Tile_X0D_Y0C_lo_out[4],Tile_X0D_Y0C_hi_out[4],Tile_X0D_Y0C_lo_out[3],Tile_X0D_Y0C_lo_out[3:2],Tile_X0D_Y0C_lo_out[2],Tile_X0D_Y0C_hi_out[2:1],Tile_X0D_Y0C_lo_out[0],Tile_X0D_Y0C_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0D_Y0C_tile_id (
    .in(Tile_X0D_Y0C_tile_id_in),
    .out(Tile_X0D_Y0C_tile_id_out)
);
Tile_PE Tile_X0D_Y0D (
    .SB_T0_EAST_SB_IN_B1(Tile_X0E_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0E_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0D_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0D_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0D_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0D_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0D_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0D_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0D_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0D_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0D_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0D_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0C_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0C_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0D_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0D_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0E_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0E_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0D_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0D_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0D_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0D_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0D_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0D_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0D_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0D_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0D_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0D_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0C_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0C_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0D_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0D_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0E_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0E_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0D_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0D_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0D_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0D_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0D_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0D_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0D_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0D_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0D_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0D_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0C_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0C_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0D_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0D_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0E_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0E_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0D_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0D_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0D_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0D_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0D_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0D_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0D_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0D_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0D_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0D_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0C_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0C_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0D_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0D_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0E_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0E_Y0D_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0D_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0D_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0D_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0D_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0D_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0D_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0D_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0D_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0D_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0D_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0C_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0C_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0D_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0D_Y0D_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0D_Y0C_clk_out),
    .clk_out(Tile_X0D_Y0D_clk_out),
    .clk_pass_through(Tile_X0D_Y0C_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0D_Y0D_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0D_Y0D_clk_pass_through_out_right),
    .config_config_addr(Tile_X0D_Y0C_config_out_config_addr),
    .config_config_data(Tile_X0D_Y0C_config_out_config_data),
    .config_out_config_addr(Tile_X0D_Y0D_config_out_config_addr),
    .config_out_config_data(Tile_X0D_Y0D_config_out_config_data),
    .config_out_read(Tile_X0D_Y0D_config_out_read),
    .config_out_write(Tile_X0D_Y0D_config_out_write),
    .config_read(Tile_X0D_Y0C_config_out_read),
    .config_write(Tile_X0D_Y0C_config_out_write),
    .hi(Tile_X0D_Y0D_hi_unq1),
    .lo(Tile_X0D_Y0D_lo_unq1),
    .read_config_data(Tile_X0D_Y0D_read_config_data),
    .read_config_data_in(Tile_X0D_Y0C_read_config_data),
    .reset(Tile_X0D_Y0C_reset_out),
    .reset_out(Tile_X0D_Y0D_reset_out),
    .stall(Tile_X0D_Y0C_stall_out),
    .stall_out(Tile_X0D_Y0D_stall_out),
    .tile_id(Tile_X0D_Y0D_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0D_Y0D_hi (
    .in(Tile_X0D_Y0D_hi_unq1),
    .out(Tile_X0D_Y0D_hi_out)
);
mantle_wire__typeBit8 Tile_X0D_Y0D_lo (
    .in(Tile_X0D_Y0D_lo_unq1),
    .out(Tile_X0D_Y0D_lo_out)
);
wire [15:0] Tile_X0D_Y0D_tile_id_out;
assign Tile_X0D_Y0D_tile_id_out = {Tile_X0D_Y0D_lo_out[7],Tile_X0D_Y0D_lo_out[7:6],Tile_X0D_Y0D_lo_out[6],Tile_X0D_Y0D_hi_out[6:5],Tile_X0D_Y0D_lo_out[4],Tile_X0D_Y0D_hi_out[4],Tile_X0D_Y0D_lo_out[3],Tile_X0D_Y0D_lo_out[3:2],Tile_X0D_Y0D_lo_out[2],Tile_X0D_Y0D_hi_out[2:1],Tile_X0D_Y0D_lo_out[0],Tile_X0D_Y0D_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X0D_Y0D_tile_id (
    .in(Tile_X0D_Y0D_tile_id_in),
    .out(Tile_X0D_Y0D_tile_id_out)
);
Tile_PE Tile_X0D_Y0E (
    .SB_T0_EAST_SB_IN_B1(Tile_X0E_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0E_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0D_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0D_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0D_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0D_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0D_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0D_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0D_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0D_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0D_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0D_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0C_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0C_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0D_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0D_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0E_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0E_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0D_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0D_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0D_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0D_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0D_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0D_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0D_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0D_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0D_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0D_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0C_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0C_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0D_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0D_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0E_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0E_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0D_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0D_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0D_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0D_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0D_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0D_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0D_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0D_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0D_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0D_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0C_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0C_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0D_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0D_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0E_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0E_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0D_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0D_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0D_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0D_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0D_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0D_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0D_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0D_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0D_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0D_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0C_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0C_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0D_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0D_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0E_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0E_Y0E_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0D_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0D_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0D_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0D_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0D_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0D_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0D_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0D_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0D_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0D_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0C_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0C_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0D_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0D_Y0E_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0D_Y0D_clk_out),
    .clk_out(Tile_X0D_Y0E_clk_out),
    .clk_pass_through(Tile_X0D_Y0D_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0D_Y0E_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0D_Y0E_clk_pass_through_out_right),
    .config_config_addr(Tile_X0D_Y0D_config_out_config_addr),
    .config_config_data(Tile_X0D_Y0D_config_out_config_data),
    .config_out_config_addr(Tile_X0D_Y0E_config_out_config_addr),
    .config_out_config_data(Tile_X0D_Y0E_config_out_config_data),
    .config_out_read(Tile_X0D_Y0E_config_out_read),
    .config_out_write(Tile_X0D_Y0E_config_out_write),
    .config_read(Tile_X0D_Y0D_config_out_read),
    .config_write(Tile_X0D_Y0D_config_out_write),
    .hi(Tile_X0D_Y0E_hi_unq1),
    .lo(Tile_X0D_Y0E_lo_unq1),
    .read_config_data(Tile_X0D_Y0E_read_config_data),
    .read_config_data_in(Tile_X0D_Y0D_read_config_data),
    .reset(Tile_X0D_Y0D_reset_out),
    .reset_out(Tile_X0D_Y0E_reset_out),
    .stall(Tile_X0D_Y0D_stall_out),
    .stall_out(Tile_X0D_Y0E_stall_out),
    .tile_id(Tile_X0D_Y0E_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0D_Y0E_hi (
    .in(Tile_X0D_Y0E_hi_unq1),
    .out(Tile_X0D_Y0E_hi_out)
);
mantle_wire__typeBit8 Tile_X0D_Y0E_lo (
    .in(Tile_X0D_Y0E_lo_unq1),
    .out(Tile_X0D_Y0E_lo_out)
);
wire [15:0] Tile_X0D_Y0E_tile_id_out;
assign Tile_X0D_Y0E_tile_id_out = {Tile_X0D_Y0E_lo_out[7],Tile_X0D_Y0E_lo_out[7:6],Tile_X0D_Y0E_lo_out[6],Tile_X0D_Y0E_hi_out[6:5],Tile_X0D_Y0E_lo_out[4],Tile_X0D_Y0E_hi_out[4],Tile_X0D_Y0E_lo_out[3],Tile_X0D_Y0E_lo_out[3:2],Tile_X0D_Y0E_lo_out[2],Tile_X0D_Y0E_hi_out[2:1],Tile_X0D_Y0E_hi_out[1],Tile_X0D_Y0E_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0D_Y0E_tile_id (
    .in(Tile_X0D_Y0E_tile_id_in),
    .out(Tile_X0D_Y0E_tile_id_out)
);
Tile_PE Tile_X0D_Y0F (
    .SB_T0_EAST_SB_IN_B1(Tile_X0E_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0E_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0D_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0D_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0D_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0D_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0D_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0D_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0D_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0D_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0D_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0D_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0C_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0C_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0D_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0D_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0E_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0E_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0D_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0D_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0D_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0D_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0D_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0D_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0D_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0D_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0D_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0D_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0C_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0C_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0D_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0D_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0E_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0E_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0D_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0D_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0D_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0D_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0D_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0D_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0D_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0D_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0D_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0D_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0C_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0C_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0D_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0D_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0E_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0E_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0D_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0D_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0D_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0D_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0D_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0D_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0D_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0D_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0D_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0D_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0C_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0C_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0D_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0D_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0E_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0E_Y0F_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0D_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0D_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0D_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0D_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0D_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0D_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0D_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0D_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0D_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0D_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0C_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0C_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0D_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0D_Y0F_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0D_Y0E_clk_out),
    .clk_out(Tile_X0D_Y0F_clk_out),
    .clk_pass_through(Tile_X0D_Y0E_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0D_Y0F_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0D_Y0F_clk_pass_through_out_right),
    .config_config_addr(Tile_X0D_Y0E_config_out_config_addr),
    .config_config_data(Tile_X0D_Y0E_config_out_config_data),
    .config_out_config_addr(Tile_X0D_Y0F_config_out_config_addr),
    .config_out_config_data(Tile_X0D_Y0F_config_out_config_data),
    .config_out_read(Tile_X0D_Y0F_config_out_read),
    .config_out_write(Tile_X0D_Y0F_config_out_write),
    .config_read(Tile_X0D_Y0E_config_out_read),
    .config_write(Tile_X0D_Y0E_config_out_write),
    .hi(Tile_X0D_Y0F_hi_unq1),
    .lo(Tile_X0D_Y0F_lo_unq1),
    .read_config_data(Tile_X0D_Y0F_read_config_data),
    .read_config_data_in(Tile_X0D_Y0E_read_config_data),
    .reset(Tile_X0D_Y0E_reset_out),
    .reset_out(Tile_X0D_Y0F_reset_out),
    .stall(Tile_X0D_Y0E_stall_out),
    .stall_out(Tile_X0D_Y0F_stall_out),
    .tile_id(Tile_X0D_Y0F_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0D_Y0F_hi (
    .in(Tile_X0D_Y0F_hi_unq1),
    .out(Tile_X0D_Y0F_hi_out)
);
mantle_wire__typeBit8 Tile_X0D_Y0F_lo (
    .in(Tile_X0D_Y0F_lo_unq1),
    .out(Tile_X0D_Y0F_lo_out)
);
wire [15:0] Tile_X0D_Y0F_tile_id_out;
assign Tile_X0D_Y0F_tile_id_out = {Tile_X0D_Y0F_lo_out[7],Tile_X0D_Y0F_lo_out[7:6],Tile_X0D_Y0F_lo_out[6],Tile_X0D_Y0F_hi_out[6:5],Tile_X0D_Y0F_lo_out[4],Tile_X0D_Y0F_hi_out[4],Tile_X0D_Y0F_lo_out[3],Tile_X0D_Y0F_lo_out[3:2],Tile_X0D_Y0F_lo_out[2],Tile_X0D_Y0F_hi_out[2:1],Tile_X0D_Y0F_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X0D_Y0F_tile_id (
    .in(Tile_X0D_Y0F_tile_id_in),
    .out(Tile_X0D_Y0F_tile_id_out)
);
Tile_PE Tile_X0D_Y10 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0E_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0E_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0D_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0D_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0D_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0D_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0D_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0D_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T0_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0D_Y10_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0D_Y10_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0C_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0C_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0D_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0D_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0E_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0E_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0D_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0D_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0D_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0D_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0D_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0D_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T1_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0D_Y10_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0D_Y10_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0C_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0C_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0D_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0D_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0E_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0E_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0D_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0D_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0D_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0D_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0D_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0D_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T2_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0D_Y10_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0D_Y10_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0C_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0C_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0D_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0D_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0E_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0E_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0D_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0D_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0D_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0D_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0D_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0D_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T3_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0D_Y10_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0D_Y10_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0C_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0C_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0D_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0D_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0E_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0E_Y10_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0D_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0D_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0D_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0D_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0D_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0D_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T4_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0D_Y10_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0D_Y10_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0C_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0C_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0D_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0D_Y10_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0D_Y0F_clk_out),
    .clk_out(Tile_X0D_Y10_clk_out),
    .clk_pass_through(Tile_X0D_Y0F_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0D_Y10_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0D_Y10_clk_pass_through_out_right),
    .config_config_addr(Tile_X0D_Y0F_config_out_config_addr),
    .config_config_data(Tile_X0D_Y0F_config_out_config_data),
    .config_out_config_addr(Tile_X0D_Y10_config_out_config_addr),
    .config_out_config_data(Tile_X0D_Y10_config_out_config_data),
    .config_out_read(Tile_X0D_Y10_config_out_read),
    .config_out_write(Tile_X0D_Y10_config_out_write),
    .config_read(Tile_X0D_Y0F_config_out_read),
    .config_write(Tile_X0D_Y0F_config_out_write),
    .hi(Tile_X0D_Y10_hi_unq1),
    .lo(Tile_X0D_Y10_lo_unq1),
    .read_config_data(Tile_X0D_Y10_read_config_data),
    .read_config_data_in(Tile_X0D_Y0F_read_config_data),
    .reset(Tile_X0D_Y0F_reset_out),
    .reset_out(Tile_X0D_Y10_reset_out),
    .stall(Tile_X0D_Y0F_stall_out),
    .stall_out(Tile_X0D_Y10_stall_out),
    .tile_id(Tile_X0D_Y10_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0D_Y10_hi (
    .in(Tile_X0D_Y10_hi_unq1),
    .out(Tile_X0D_Y10_hi_out)
);
mantle_wire__typeBit8 Tile_X0D_Y10_lo (
    .in(Tile_X0D_Y10_lo_unq1),
    .out(Tile_X0D_Y10_lo_out)
);
wire [15:0] Tile_X0D_Y10_tile_id_out;
assign Tile_X0D_Y10_tile_id_out = {Tile_X0D_Y10_lo_out[7],Tile_X0D_Y10_lo_out[7:6],Tile_X0D_Y10_lo_out[6],Tile_X0D_Y10_hi_out[6:5],Tile_X0D_Y10_lo_out[4],Tile_X0D_Y10_hi_out[4],Tile_X0D_Y10_lo_out[3],Tile_X0D_Y10_lo_out[3:2],Tile_X0D_Y10_hi_out[2],Tile_X0D_Y10_lo_out[1],Tile_X0D_Y10_lo_out[1:0],Tile_X0D_Y10_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0D_Y10_tile_id (
    .in(Tile_X0D_Y10_tile_id_in),
    .out(Tile_X0D_Y10_tile_id_out)
);
wire [15:0] Tile_X0E_Y00_tile_id;
assign Tile_X0E_Y00_tile_id = {Tile_X0E_Y00_lo[7],Tile_X0E_Y00_lo[7:6],Tile_X0E_Y00_lo[6],Tile_X0E_Y00_hi[6:5],Tile_X0E_Y00_hi[5],Tile_X0E_Y00_lo[4:3],Tile_X0E_Y00_lo[3:2],Tile_X0E_Y00_lo[2:1],Tile_X0E_Y00_lo[1:0],Tile_X0E_Y00_lo[0]};
Tile_io_core Tile_X0E_Y00 (
    .tile_id(Tile_X0E_Y00_tile_id),
    .glb2io_1(glb2io_1_X0E_Y00),
    .f2io_1(Tile_X0E_Y01_SB_T0_NORTH_SB_OUT_B1),
    .io2glb_1(Tile_X0E_Y00_io2glb_1),
    .io2f_1(Tile_X0E_Y00_io2f_1),
    .glb2io_16(glb2io_16_X0E_Y00),
    .f2io_16(Tile_X0E_Y01_SB_T0_NORTH_SB_OUT_B16),
    .io2glb_16(Tile_X0E_Y00_io2glb_16),
    .io2f_16(Tile_X0E_Y00_io2f_16),
    .hi(Tile_X0E_Y00_hi),
    .lo(Tile_X0E_Y00_lo)
);
Tile_PE Tile_X0E_Y01 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0F_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0F_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0E_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0E_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0E_Y00_io2f_1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0E_Y00_io2f_16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0E_Y01_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0E_Y01_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0E_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0E_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0E_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0E_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0D_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0D_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0E_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0E_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0F_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0F_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0E_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0E_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0E_Y00_io2f_1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0E_Y00_io2f_16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0E_Y01_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0E_Y01_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0E_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0E_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0E_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0E_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0D_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0D_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0E_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0E_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0F_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0F_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0E_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0E_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0E_Y00_io2f_1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0E_Y00_io2f_16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0E_Y01_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0E_Y01_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0E_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0E_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0E_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0E_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0D_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0D_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0E_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0E_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0F_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0F_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0E_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0E_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0E_Y00_io2f_1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0E_Y00_io2f_16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0E_Y01_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0E_Y01_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0E_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0E_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0E_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0E_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0D_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0D_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0E_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0E_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0F_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0F_Y01_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0E_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0E_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0E_Y00_io2f_1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0E_Y00_io2f_16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0E_Y01_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0E_Y01_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0E_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0E_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0E_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0E_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0D_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0D_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0E_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0E_Y01_SB_T4_WEST_SB_OUT_B16),
    .clk(clk),
    .clk_out(Tile_X0E_Y01_clk_out),
    .clk_pass_through(clk),
    .clk_pass_through_out_bot(Tile_X0E_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0E_Y01_clk_pass_through_out_right),
    .config_config_addr(config_14_config_addr),
    .config_config_data(config_14_config_data),
    .config_out_config_addr(Tile_X0E_Y01_config_out_config_addr),
    .config_out_config_data(Tile_X0E_Y01_config_out_config_data),
    .config_out_read(Tile_X0E_Y01_config_out_read),
    .config_out_write(Tile_X0E_Y01_config_out_write),
    .config_read(config_14_read),
    .config_write(config_14_write),
    .hi(Tile_X0E_Y01_hi_unq1),
    .lo(Tile_X0E_Y01_lo_unq1),
    .read_config_data(Tile_X0E_Y01_read_config_data),
    .read_config_data_in(const_0_32_out),
    .reset(reset),
    .reset_out(Tile_X0E_Y01_reset_out),
    .stall(stall[14]),
    .stall_out(Tile_X0E_Y01_stall_out),
    .tile_id(Tile_X0E_Y01_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0E_Y01_hi (
    .in(Tile_X0E_Y01_hi_unq1),
    .out(Tile_X0E_Y01_hi_out)
);
mantle_wire__typeBit8 Tile_X0E_Y01_lo (
    .in(Tile_X0E_Y01_lo_unq1),
    .out(Tile_X0E_Y01_lo_out)
);
wire [15:0] Tile_X0E_Y01_tile_id_out;
assign Tile_X0E_Y01_tile_id_out = {Tile_X0E_Y01_lo_out[7],Tile_X0E_Y01_lo_out[7:6],Tile_X0E_Y01_lo_out[6],Tile_X0E_Y01_hi_out[6:5],Tile_X0E_Y01_hi_out[5],Tile_X0E_Y01_lo_out[4:3],Tile_X0E_Y01_lo_out[3:2],Tile_X0E_Y01_lo_out[2:1],Tile_X0E_Y01_lo_out[1:0],Tile_X0E_Y01_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X0E_Y01_tile_id (
    .in(Tile_X0E_Y01_tile_id_in),
    .out(Tile_X0E_Y01_tile_id_out)
);
Tile_PE Tile_X0E_Y02 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0F_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0F_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0E_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0E_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0E_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0E_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0E_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0E_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0E_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0E_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0E_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0E_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0D_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0D_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0E_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0E_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0F_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0F_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0E_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0E_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0E_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0E_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0E_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0E_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0E_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0E_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0E_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0E_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0D_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0D_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0E_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0E_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0F_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0F_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0E_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0E_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0E_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0E_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0E_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0E_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0E_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0E_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0E_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0E_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0D_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0D_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0E_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0E_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0F_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0F_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0E_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0E_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0E_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0E_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0E_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0E_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0E_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0E_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0E_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0E_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0D_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0D_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0E_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0E_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0F_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0F_Y02_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0E_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0E_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0E_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0E_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0E_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0E_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0E_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0E_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0E_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0E_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0D_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0D_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0E_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0E_Y02_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y01_clk_out),
    .clk_out(Tile_X0E_Y02_clk_out),
    .clk_pass_through(Tile_X0E_Y01_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0E_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0E_Y02_clk_pass_through_out_right),
    .config_config_addr(Tile_X0E_Y01_config_out_config_addr),
    .config_config_data(Tile_X0E_Y01_config_out_config_data),
    .config_out_config_addr(Tile_X0E_Y02_config_out_config_addr),
    .config_out_config_data(Tile_X0E_Y02_config_out_config_data),
    .config_out_read(Tile_X0E_Y02_config_out_read),
    .config_out_write(Tile_X0E_Y02_config_out_write),
    .config_read(Tile_X0E_Y01_config_out_read),
    .config_write(Tile_X0E_Y01_config_out_write),
    .hi(Tile_X0E_Y02_hi_unq1),
    .lo(Tile_X0E_Y02_lo_unq1),
    .read_config_data(Tile_X0E_Y02_read_config_data),
    .read_config_data_in(Tile_X0E_Y01_read_config_data),
    .reset(Tile_X0E_Y01_reset_out),
    .reset_out(Tile_X0E_Y02_reset_out),
    .stall(Tile_X0E_Y01_stall_out),
    .stall_out(Tile_X0E_Y02_stall_out),
    .tile_id(Tile_X0E_Y02_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0E_Y02_hi (
    .in(Tile_X0E_Y02_hi_unq1),
    .out(Tile_X0E_Y02_hi_out)
);
mantle_wire__typeBit8 Tile_X0E_Y02_lo (
    .in(Tile_X0E_Y02_lo_unq1),
    .out(Tile_X0E_Y02_lo_out)
);
wire [15:0] Tile_X0E_Y02_tile_id_out;
assign Tile_X0E_Y02_tile_id_out = {Tile_X0E_Y02_lo_out[7],Tile_X0E_Y02_lo_out[7:6],Tile_X0E_Y02_lo_out[6],Tile_X0E_Y02_hi_out[6:5],Tile_X0E_Y02_hi_out[5],Tile_X0E_Y02_lo_out[4:3],Tile_X0E_Y02_lo_out[3:2],Tile_X0E_Y02_lo_out[2:1],Tile_X0E_Y02_lo_out[1],Tile_X0E_Y02_hi_out[1],Tile_X0E_Y02_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0E_Y02_tile_id (
    .in(Tile_X0E_Y02_tile_id_in),
    .out(Tile_X0E_Y02_tile_id_out)
);
Tile_PE Tile_X0E_Y03 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0F_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0F_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0E_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0E_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0E_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0E_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0E_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0E_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0E_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0E_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0E_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0E_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0D_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0D_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0E_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0E_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0F_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0F_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0E_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0E_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0E_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0E_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0E_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0E_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0E_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0E_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0E_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0E_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0D_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0D_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0E_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0E_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0F_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0F_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0E_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0E_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0E_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0E_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0E_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0E_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0E_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0E_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0E_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0E_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0D_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0D_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0E_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0E_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0F_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0F_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0E_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0E_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0E_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0E_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0E_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0E_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0E_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0E_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0E_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0E_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0D_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0D_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0E_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0E_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0F_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0F_Y03_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0E_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0E_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0E_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0E_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0E_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0E_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0E_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0E_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0E_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0E_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0D_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0D_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0E_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0E_Y03_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y02_clk_out),
    .clk_out(Tile_X0E_Y03_clk_out),
    .clk_pass_through(Tile_X0E_Y02_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0E_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0E_Y03_clk_pass_through_out_right),
    .config_config_addr(Tile_X0E_Y02_config_out_config_addr),
    .config_config_data(Tile_X0E_Y02_config_out_config_data),
    .config_out_config_addr(Tile_X0E_Y03_config_out_config_addr),
    .config_out_config_data(Tile_X0E_Y03_config_out_config_data),
    .config_out_read(Tile_X0E_Y03_config_out_read),
    .config_out_write(Tile_X0E_Y03_config_out_write),
    .config_read(Tile_X0E_Y02_config_out_read),
    .config_write(Tile_X0E_Y02_config_out_write),
    .hi(Tile_X0E_Y03_hi_unq1),
    .lo(Tile_X0E_Y03_lo_unq1),
    .read_config_data(Tile_X0E_Y03_read_config_data),
    .read_config_data_in(Tile_X0E_Y02_read_config_data),
    .reset(Tile_X0E_Y02_reset_out),
    .reset_out(Tile_X0E_Y03_reset_out),
    .stall(Tile_X0E_Y02_stall_out),
    .stall_out(Tile_X0E_Y03_stall_out),
    .tile_id(Tile_X0E_Y03_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0E_Y03_hi (
    .in(Tile_X0E_Y03_hi_unq1),
    .out(Tile_X0E_Y03_hi_out)
);
mantle_wire__typeBit8 Tile_X0E_Y03_lo (
    .in(Tile_X0E_Y03_lo_unq1),
    .out(Tile_X0E_Y03_lo_out)
);
wire [15:0] Tile_X0E_Y03_tile_id_out;
assign Tile_X0E_Y03_tile_id_out = {Tile_X0E_Y03_lo_out[7],Tile_X0E_Y03_lo_out[7:6],Tile_X0E_Y03_lo_out[6],Tile_X0E_Y03_hi_out[6:5],Tile_X0E_Y03_hi_out[5],Tile_X0E_Y03_lo_out[4:3],Tile_X0E_Y03_lo_out[3:2],Tile_X0E_Y03_lo_out[2:1],Tile_X0E_Y03_lo_out[1],Tile_X0E_Y03_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X0E_Y03_tile_id (
    .in(Tile_X0E_Y03_tile_id_in),
    .out(Tile_X0E_Y03_tile_id_out)
);
Tile_PE Tile_X0E_Y04 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0F_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0F_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0E_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0E_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0E_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0E_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0E_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0E_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0E_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0E_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0E_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0E_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0D_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0D_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0E_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0E_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0F_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0F_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0E_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0E_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0E_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0E_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0E_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0E_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0E_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0E_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0E_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0E_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0D_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0D_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0E_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0E_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0F_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0F_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0E_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0E_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0E_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0E_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0E_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0E_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0E_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0E_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0E_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0E_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0D_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0D_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0E_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0E_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0F_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0F_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0E_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0E_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0E_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0E_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0E_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0E_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0E_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0E_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0E_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0E_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0D_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0D_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0E_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0E_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0F_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0F_Y04_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0E_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0E_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0E_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0E_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0E_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0E_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0E_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0E_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0E_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0E_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0D_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0D_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0E_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0E_Y04_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y03_clk_out),
    .clk_out(Tile_X0E_Y04_clk_out),
    .clk_pass_through(Tile_X0E_Y03_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0E_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0E_Y04_clk_pass_through_out_right),
    .config_config_addr(Tile_X0E_Y03_config_out_config_addr),
    .config_config_data(Tile_X0E_Y03_config_out_config_data),
    .config_out_config_addr(Tile_X0E_Y04_config_out_config_addr),
    .config_out_config_data(Tile_X0E_Y04_config_out_config_data),
    .config_out_read(Tile_X0E_Y04_config_out_read),
    .config_out_write(Tile_X0E_Y04_config_out_write),
    .config_read(Tile_X0E_Y03_config_out_read),
    .config_write(Tile_X0E_Y03_config_out_write),
    .hi(Tile_X0E_Y04_hi_unq1),
    .lo(Tile_X0E_Y04_lo_unq1),
    .read_config_data(Tile_X0E_Y04_read_config_data),
    .read_config_data_in(Tile_X0E_Y03_read_config_data),
    .reset(Tile_X0E_Y03_reset_out),
    .reset_out(Tile_X0E_Y04_reset_out),
    .stall(Tile_X0E_Y03_stall_out),
    .stall_out(Tile_X0E_Y04_stall_out),
    .tile_id(Tile_X0E_Y04_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0E_Y04_hi (
    .in(Tile_X0E_Y04_hi_unq1),
    .out(Tile_X0E_Y04_hi_out)
);
mantle_wire__typeBit8 Tile_X0E_Y04_lo (
    .in(Tile_X0E_Y04_lo_unq1),
    .out(Tile_X0E_Y04_lo_out)
);
wire [15:0] Tile_X0E_Y04_tile_id_out;
assign Tile_X0E_Y04_tile_id_out = {Tile_X0E_Y04_lo_out[7],Tile_X0E_Y04_lo_out[7:6],Tile_X0E_Y04_lo_out[6],Tile_X0E_Y04_hi_out[6:5],Tile_X0E_Y04_hi_out[5],Tile_X0E_Y04_lo_out[4:3],Tile_X0E_Y04_lo_out[3:2],Tile_X0E_Y04_lo_out[2:1],Tile_X0E_Y04_hi_out[1],Tile_X0E_Y04_lo_out[0],Tile_X0E_Y04_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0E_Y04_tile_id (
    .in(Tile_X0E_Y04_tile_id_in),
    .out(Tile_X0E_Y04_tile_id_out)
);
Tile_PE Tile_X0E_Y05 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0F_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0F_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0E_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0E_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0E_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0E_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0E_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0E_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0E_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0E_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0E_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0E_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0D_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0D_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0E_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0E_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0F_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0F_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0E_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0E_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0E_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0E_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0E_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0E_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0E_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0E_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0E_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0E_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0D_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0D_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0E_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0E_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0F_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0F_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0E_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0E_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0E_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0E_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0E_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0E_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0E_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0E_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0E_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0E_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0D_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0D_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0E_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0E_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0F_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0F_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0E_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0E_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0E_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0E_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0E_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0E_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0E_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0E_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0E_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0E_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0D_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0D_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0E_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0E_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0F_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0F_Y05_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0E_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0E_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0E_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0E_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0E_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0E_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0E_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0E_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0E_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0E_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0D_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0D_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0E_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0E_Y05_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y04_clk_out),
    .clk_out(Tile_X0E_Y05_clk_out),
    .clk_pass_through(Tile_X0E_Y04_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0E_Y05_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0E_Y05_clk_pass_through_out_right),
    .config_config_addr(Tile_X0E_Y04_config_out_config_addr),
    .config_config_data(Tile_X0E_Y04_config_out_config_data),
    .config_out_config_addr(Tile_X0E_Y05_config_out_config_addr),
    .config_out_config_data(Tile_X0E_Y05_config_out_config_data),
    .config_out_read(Tile_X0E_Y05_config_out_read),
    .config_out_write(Tile_X0E_Y05_config_out_write),
    .config_read(Tile_X0E_Y04_config_out_read),
    .config_write(Tile_X0E_Y04_config_out_write),
    .hi(Tile_X0E_Y05_hi_unq1),
    .lo(Tile_X0E_Y05_lo_unq1),
    .read_config_data(Tile_X0E_Y05_read_config_data),
    .read_config_data_in(Tile_X0E_Y04_read_config_data),
    .reset(Tile_X0E_Y04_reset_out),
    .reset_out(Tile_X0E_Y05_reset_out),
    .stall(Tile_X0E_Y04_stall_out),
    .stall_out(Tile_X0E_Y05_stall_out),
    .tile_id(Tile_X0E_Y05_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0E_Y05_hi (
    .in(Tile_X0E_Y05_hi_unq1),
    .out(Tile_X0E_Y05_hi_out)
);
mantle_wire__typeBit8 Tile_X0E_Y05_lo (
    .in(Tile_X0E_Y05_lo_unq1),
    .out(Tile_X0E_Y05_lo_out)
);
wire [15:0] Tile_X0E_Y05_tile_id_out;
assign Tile_X0E_Y05_tile_id_out = {Tile_X0E_Y05_lo_out[7],Tile_X0E_Y05_lo_out[7:6],Tile_X0E_Y05_lo_out[6],Tile_X0E_Y05_hi_out[6:5],Tile_X0E_Y05_hi_out[5],Tile_X0E_Y05_lo_out[4:3],Tile_X0E_Y05_lo_out[3:2],Tile_X0E_Y05_lo_out[2:1],Tile_X0E_Y05_hi_out[1],Tile_X0E_Y05_lo_out[0],Tile_X0E_Y05_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X0E_Y05_tile_id (
    .in(Tile_X0E_Y05_tile_id_in),
    .out(Tile_X0E_Y05_tile_id_out)
);
Tile_PE Tile_X0E_Y06 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0F_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0F_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0E_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0E_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0E_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0E_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0E_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0E_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0E_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0E_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0E_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0E_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0D_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0D_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0E_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0E_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0F_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0F_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0E_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0E_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0E_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0E_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0E_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0E_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0E_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0E_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0E_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0E_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0D_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0D_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0E_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0E_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0F_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0F_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0E_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0E_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0E_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0E_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0E_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0E_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0E_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0E_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0E_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0E_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0D_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0D_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0E_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0E_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0F_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0F_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0E_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0E_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0E_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0E_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0E_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0E_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0E_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0E_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0E_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0E_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0D_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0D_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0E_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0E_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0F_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0F_Y06_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0E_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0E_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0E_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0E_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0E_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0E_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0E_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0E_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0E_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0E_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0D_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0D_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0E_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0E_Y06_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y05_clk_out),
    .clk_out(Tile_X0E_Y06_clk_out),
    .clk_pass_through(Tile_X0E_Y05_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0E_Y06_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0E_Y06_clk_pass_through_out_right),
    .config_config_addr(Tile_X0E_Y05_config_out_config_addr),
    .config_config_data(Tile_X0E_Y05_config_out_config_data),
    .config_out_config_addr(Tile_X0E_Y06_config_out_config_addr),
    .config_out_config_data(Tile_X0E_Y06_config_out_config_data),
    .config_out_read(Tile_X0E_Y06_config_out_read),
    .config_out_write(Tile_X0E_Y06_config_out_write),
    .config_read(Tile_X0E_Y05_config_out_read),
    .config_write(Tile_X0E_Y05_config_out_write),
    .hi(Tile_X0E_Y06_hi_unq1),
    .lo(Tile_X0E_Y06_lo_unq1),
    .read_config_data(Tile_X0E_Y06_read_config_data),
    .read_config_data_in(Tile_X0E_Y05_read_config_data),
    .reset(Tile_X0E_Y05_reset_out),
    .reset_out(Tile_X0E_Y06_reset_out),
    .stall(Tile_X0E_Y05_stall_out),
    .stall_out(Tile_X0E_Y06_stall_out),
    .tile_id(Tile_X0E_Y06_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0E_Y06_hi (
    .in(Tile_X0E_Y06_hi_unq1),
    .out(Tile_X0E_Y06_hi_out)
);
mantle_wire__typeBit8 Tile_X0E_Y06_lo (
    .in(Tile_X0E_Y06_lo_unq1),
    .out(Tile_X0E_Y06_lo_out)
);
wire [15:0] Tile_X0E_Y06_tile_id_out;
assign Tile_X0E_Y06_tile_id_out = {Tile_X0E_Y06_lo_out[7],Tile_X0E_Y06_lo_out[7:6],Tile_X0E_Y06_lo_out[6],Tile_X0E_Y06_hi_out[6:5],Tile_X0E_Y06_hi_out[5],Tile_X0E_Y06_lo_out[4:3],Tile_X0E_Y06_lo_out[3:2],Tile_X0E_Y06_lo_out[2:1],Tile_X0E_Y06_hi_out[1],Tile_X0E_Y06_hi_out[1],Tile_X0E_Y06_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0E_Y06_tile_id (
    .in(Tile_X0E_Y06_tile_id_in),
    .out(Tile_X0E_Y06_tile_id_out)
);
Tile_PE Tile_X0E_Y07 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0F_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0F_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0E_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0E_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0E_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0E_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0E_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0E_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0E_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0E_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0E_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0E_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0D_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0D_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0E_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0E_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0F_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0F_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0E_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0E_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0E_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0E_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0E_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0E_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0E_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0E_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0E_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0E_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0D_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0D_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0E_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0E_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0F_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0F_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0E_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0E_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0E_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0E_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0E_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0E_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0E_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0E_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0E_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0E_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0D_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0D_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0E_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0E_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0F_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0F_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0E_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0E_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0E_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0E_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0E_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0E_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0E_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0E_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0E_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0E_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0D_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0D_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0E_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0E_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0F_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0F_Y07_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0E_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0E_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0E_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0E_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0E_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0E_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0E_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0E_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0E_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0E_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0D_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0D_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0E_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0E_Y07_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y06_clk_out),
    .clk_out(Tile_X0E_Y07_clk_out),
    .clk_pass_through(Tile_X0E_Y06_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0E_Y07_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0E_Y07_clk_pass_through_out_right),
    .config_config_addr(Tile_X0E_Y06_config_out_config_addr),
    .config_config_data(Tile_X0E_Y06_config_out_config_data),
    .config_out_config_addr(Tile_X0E_Y07_config_out_config_addr),
    .config_out_config_data(Tile_X0E_Y07_config_out_config_data),
    .config_out_read(Tile_X0E_Y07_config_out_read),
    .config_out_write(Tile_X0E_Y07_config_out_write),
    .config_read(Tile_X0E_Y06_config_out_read),
    .config_write(Tile_X0E_Y06_config_out_write),
    .hi(Tile_X0E_Y07_hi_unq1),
    .lo(Tile_X0E_Y07_lo_unq1),
    .read_config_data(Tile_X0E_Y07_read_config_data),
    .read_config_data_in(Tile_X0E_Y06_read_config_data),
    .reset(Tile_X0E_Y06_reset_out),
    .reset_out(Tile_X0E_Y07_reset_out),
    .stall(Tile_X0E_Y06_stall_out),
    .stall_out(Tile_X0E_Y07_stall_out),
    .tile_id(Tile_X0E_Y07_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0E_Y07_hi (
    .in(Tile_X0E_Y07_hi_unq1),
    .out(Tile_X0E_Y07_hi_out)
);
mantle_wire__typeBit8 Tile_X0E_Y07_lo (
    .in(Tile_X0E_Y07_lo_unq1),
    .out(Tile_X0E_Y07_lo_out)
);
wire [15:0] Tile_X0E_Y07_tile_id_out;
assign Tile_X0E_Y07_tile_id_out = {Tile_X0E_Y07_lo_out[7],Tile_X0E_Y07_lo_out[7:6],Tile_X0E_Y07_lo_out[6],Tile_X0E_Y07_hi_out[6:5],Tile_X0E_Y07_hi_out[5],Tile_X0E_Y07_lo_out[4:3],Tile_X0E_Y07_lo_out[3:2],Tile_X0E_Y07_lo_out[2:1],Tile_X0E_Y07_hi_out[1],Tile_X0E_Y07_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X0E_Y07_tile_id (
    .in(Tile_X0E_Y07_tile_id_in),
    .out(Tile_X0E_Y07_tile_id_out)
);
Tile_PE Tile_X0E_Y08 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0F_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0F_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0E_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0E_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0E_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0E_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0E_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0E_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0E_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0E_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0E_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0E_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0D_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0D_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0E_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0E_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0F_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0F_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0E_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0E_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0E_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0E_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0E_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0E_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0E_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0E_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0E_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0E_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0D_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0D_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0E_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0E_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0F_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0F_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0E_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0E_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0E_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0E_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0E_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0E_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0E_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0E_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0E_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0E_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0D_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0D_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0E_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0E_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0F_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0F_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0E_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0E_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0E_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0E_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0E_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0E_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0E_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0E_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0E_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0E_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0D_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0D_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0E_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0E_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0F_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0F_Y08_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0E_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0E_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0E_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0E_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0E_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0E_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0E_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0E_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0E_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0E_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0D_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0D_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0E_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0E_Y08_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y07_clk_out),
    .clk_out(Tile_X0E_Y08_clk_out),
    .clk_pass_through(Tile_X0E_Y07_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0E_Y08_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0E_Y08_clk_pass_through_out_right),
    .config_config_addr(Tile_X0E_Y07_config_out_config_addr),
    .config_config_data(Tile_X0E_Y07_config_out_config_data),
    .config_out_config_addr(Tile_X0E_Y08_config_out_config_addr),
    .config_out_config_data(Tile_X0E_Y08_config_out_config_data),
    .config_out_read(Tile_X0E_Y08_config_out_read),
    .config_out_write(Tile_X0E_Y08_config_out_write),
    .config_read(Tile_X0E_Y07_config_out_read),
    .config_write(Tile_X0E_Y07_config_out_write),
    .hi(Tile_X0E_Y08_hi_unq1),
    .lo(Tile_X0E_Y08_lo_unq1),
    .read_config_data(Tile_X0E_Y08_read_config_data),
    .read_config_data_in(Tile_X0E_Y07_read_config_data),
    .reset(Tile_X0E_Y07_reset_out),
    .reset_out(Tile_X0E_Y08_reset_out),
    .stall(Tile_X0E_Y07_stall_out),
    .stall_out(Tile_X0E_Y08_stall_out),
    .tile_id(Tile_X0E_Y08_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0E_Y08_hi (
    .in(Tile_X0E_Y08_hi_unq1),
    .out(Tile_X0E_Y08_hi_out)
);
mantle_wire__typeBit8 Tile_X0E_Y08_lo (
    .in(Tile_X0E_Y08_lo_unq1),
    .out(Tile_X0E_Y08_lo_out)
);
wire [15:0] Tile_X0E_Y08_tile_id_out;
assign Tile_X0E_Y08_tile_id_out = {Tile_X0E_Y08_lo_out[7],Tile_X0E_Y08_lo_out[7:6],Tile_X0E_Y08_lo_out[6],Tile_X0E_Y08_hi_out[6:5],Tile_X0E_Y08_hi_out[5],Tile_X0E_Y08_lo_out[4:3],Tile_X0E_Y08_lo_out[3:2],Tile_X0E_Y08_lo_out[2],Tile_X0E_Y08_hi_out[2],Tile_X0E_Y08_lo_out[1:0],Tile_X0E_Y08_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0E_Y08_tile_id (
    .in(Tile_X0E_Y08_tile_id_in),
    .out(Tile_X0E_Y08_tile_id_out)
);
Tile_PE Tile_X0E_Y09 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0F_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0F_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0E_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0E_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0E_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0E_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0E_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0E_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0E_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0E_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0E_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0E_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0D_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0D_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0E_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0E_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0F_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0F_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0E_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0E_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0E_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0E_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0E_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0E_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0E_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0E_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0E_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0E_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0D_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0D_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0E_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0E_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0F_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0F_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0E_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0E_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0E_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0E_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0E_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0E_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0E_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0E_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0E_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0E_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0D_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0D_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0E_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0E_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0F_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0F_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0E_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0E_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0E_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0E_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0E_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0E_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0E_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0E_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0E_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0E_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0D_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0D_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0E_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0E_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0F_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0F_Y09_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0E_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0E_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0E_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0E_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0E_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0E_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0E_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0E_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0E_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0E_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0D_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0D_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0E_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0E_Y09_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y08_clk_out),
    .clk_out(Tile_X0E_Y09_clk_out),
    .clk_pass_through(Tile_X0E_Y08_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0E_Y09_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0E_Y09_clk_pass_through_out_right),
    .config_config_addr(ConfigPipeStage_inst14_config_out_config_addr),
    .config_config_data(ConfigPipeStage_inst14_config_out_config_data),
    .config_out_config_addr(Tile_X0E_Y09_config_out_config_addr),
    .config_out_config_data(Tile_X0E_Y09_config_out_config_data),
    .config_out_read(Tile_X0E_Y09_config_out_read),
    .config_out_write(Tile_X0E_Y09_config_out_write),
    .config_read(ConfigPipeStage_inst14_config_out_read),
    .config_write(ConfigPipeStage_inst14_config_out_write),
    .hi(Tile_X0E_Y09_hi_unq1),
    .lo(Tile_X0E_Y09_lo_unq1),
    .read_config_data(Tile_X0E_Y09_read_config_data),
    .read_config_data_in(Tile_X0E_Y08_read_config_data),
    .reset(Tile_X0E_Y08_reset_out),
    .reset_out(Tile_X0E_Y09_reset_out),
    .stall(Tile_X0E_Y08_stall_out),
    .stall_out(Tile_X0E_Y09_stall_out),
    .tile_id(Tile_X0E_Y09_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0E_Y09_hi (
    .in(Tile_X0E_Y09_hi_unq1),
    .out(Tile_X0E_Y09_hi_out)
);
mantle_wire__typeBit8 Tile_X0E_Y09_lo (
    .in(Tile_X0E_Y09_lo_unq1),
    .out(Tile_X0E_Y09_lo_out)
);
wire [15:0] Tile_X0E_Y09_tile_id_out;
assign Tile_X0E_Y09_tile_id_out = {Tile_X0E_Y09_lo_out[7],Tile_X0E_Y09_lo_out[7:6],Tile_X0E_Y09_lo_out[6],Tile_X0E_Y09_hi_out[6:5],Tile_X0E_Y09_hi_out[5],Tile_X0E_Y09_lo_out[4:3],Tile_X0E_Y09_lo_out[3:2],Tile_X0E_Y09_lo_out[2],Tile_X0E_Y09_hi_out[2],Tile_X0E_Y09_lo_out[1:0],Tile_X0E_Y09_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X0E_Y09_tile_id (
    .in(Tile_X0E_Y09_tile_id_in),
    .out(Tile_X0E_Y09_tile_id_out)
);
Tile_PE Tile_X0E_Y0A (
    .SB_T0_EAST_SB_IN_B1(Tile_X0F_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0F_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0E_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0E_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0E_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0E_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0E_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0E_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0E_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0E_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0E_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0E_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0D_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0D_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0E_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0E_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0F_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0F_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0E_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0E_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0E_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0E_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0E_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0E_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0E_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0E_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0E_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0E_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0D_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0D_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0E_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0E_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0F_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0F_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0E_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0E_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0E_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0E_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0E_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0E_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0E_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0E_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0E_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0E_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0D_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0D_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0E_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0E_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0F_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0F_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0E_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0E_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0E_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0E_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0E_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0E_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0E_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0E_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0E_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0E_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0D_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0D_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0E_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0E_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0F_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0F_Y0A_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0E_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0E_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0E_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0E_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0E_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0E_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0E_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0E_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0E_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0E_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0D_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0D_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0E_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0E_Y0A_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y09_clk_out),
    .clk_out(Tile_X0E_Y0A_clk_out),
    .clk_pass_through(Tile_X0E_Y09_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0E_Y0A_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0E_Y0A_clk_pass_through_out_right),
    .config_config_addr(Tile_X0E_Y09_config_out_config_addr),
    .config_config_data(Tile_X0E_Y09_config_out_config_data),
    .config_out_config_addr(Tile_X0E_Y0A_config_out_config_addr),
    .config_out_config_data(Tile_X0E_Y0A_config_out_config_data),
    .config_out_read(Tile_X0E_Y0A_config_out_read),
    .config_out_write(Tile_X0E_Y0A_config_out_write),
    .config_read(Tile_X0E_Y09_config_out_read),
    .config_write(Tile_X0E_Y09_config_out_write),
    .hi(Tile_X0E_Y0A_hi_unq1),
    .lo(Tile_X0E_Y0A_lo_unq1),
    .read_config_data(Tile_X0E_Y0A_read_config_data),
    .read_config_data_in(Tile_X0E_Y09_read_config_data),
    .reset(Tile_X0E_Y09_reset_out),
    .reset_out(Tile_X0E_Y0A_reset_out),
    .stall(Tile_X0E_Y09_stall_out),
    .stall_out(Tile_X0E_Y0A_stall_out),
    .tile_id(Tile_X0E_Y0A_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0E_Y0A_hi (
    .in(Tile_X0E_Y0A_hi_unq1),
    .out(Tile_X0E_Y0A_hi_out)
);
mantle_wire__typeBit8 Tile_X0E_Y0A_lo (
    .in(Tile_X0E_Y0A_lo_unq1),
    .out(Tile_X0E_Y0A_lo_out)
);
wire [15:0] Tile_X0E_Y0A_tile_id_out;
assign Tile_X0E_Y0A_tile_id_out = {Tile_X0E_Y0A_lo_out[7],Tile_X0E_Y0A_lo_out[7:6],Tile_X0E_Y0A_lo_out[6],Tile_X0E_Y0A_hi_out[6:5],Tile_X0E_Y0A_hi_out[5],Tile_X0E_Y0A_lo_out[4:3],Tile_X0E_Y0A_lo_out[3:2],Tile_X0E_Y0A_lo_out[2],Tile_X0E_Y0A_hi_out[2],Tile_X0E_Y0A_lo_out[1],Tile_X0E_Y0A_hi_out[1],Tile_X0E_Y0A_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0E_Y0A_tile_id (
    .in(Tile_X0E_Y0A_tile_id_in),
    .out(Tile_X0E_Y0A_tile_id_out)
);
Tile_PE Tile_X0E_Y0B (
    .SB_T0_EAST_SB_IN_B1(Tile_X0F_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0F_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0E_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0E_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0E_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0E_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0E_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0E_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0E_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0E_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0E_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0E_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0D_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0D_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0E_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0E_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0F_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0F_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0E_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0E_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0E_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0E_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0E_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0E_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0E_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0E_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0E_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0E_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0D_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0D_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0E_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0E_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0F_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0F_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0E_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0E_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0E_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0E_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0E_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0E_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0E_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0E_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0E_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0E_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0D_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0D_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0E_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0E_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0F_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0F_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0E_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0E_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0E_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0E_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0E_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0E_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0E_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0E_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0E_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0E_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0D_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0D_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0E_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0E_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0F_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0F_Y0B_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0E_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0E_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0E_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0E_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0E_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0E_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0E_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0E_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0E_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0E_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0D_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0D_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0E_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0E_Y0B_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y0A_clk_out),
    .clk_out(Tile_X0E_Y0B_clk_out),
    .clk_pass_through(Tile_X0E_Y0A_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0E_Y0B_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0E_Y0B_clk_pass_through_out_right),
    .config_config_addr(Tile_X0E_Y0A_config_out_config_addr),
    .config_config_data(Tile_X0E_Y0A_config_out_config_data),
    .config_out_config_addr(Tile_X0E_Y0B_config_out_config_addr),
    .config_out_config_data(Tile_X0E_Y0B_config_out_config_data),
    .config_out_read(Tile_X0E_Y0B_config_out_read),
    .config_out_write(Tile_X0E_Y0B_config_out_write),
    .config_read(Tile_X0E_Y0A_config_out_read),
    .config_write(Tile_X0E_Y0A_config_out_write),
    .hi(Tile_X0E_Y0B_hi_unq1),
    .lo(Tile_X0E_Y0B_lo_unq1),
    .read_config_data(Tile_X0E_Y0B_read_config_data),
    .read_config_data_in(Tile_X0E_Y0A_read_config_data),
    .reset(Tile_X0E_Y0A_reset_out),
    .reset_out(Tile_X0E_Y0B_reset_out),
    .stall(Tile_X0E_Y0A_stall_out),
    .stall_out(Tile_X0E_Y0B_stall_out),
    .tile_id(Tile_X0E_Y0B_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0E_Y0B_hi (
    .in(Tile_X0E_Y0B_hi_unq1),
    .out(Tile_X0E_Y0B_hi_out)
);
mantle_wire__typeBit8 Tile_X0E_Y0B_lo (
    .in(Tile_X0E_Y0B_lo_unq1),
    .out(Tile_X0E_Y0B_lo_out)
);
wire [15:0] Tile_X0E_Y0B_tile_id_out;
assign Tile_X0E_Y0B_tile_id_out = {Tile_X0E_Y0B_lo_out[7],Tile_X0E_Y0B_lo_out[7:6],Tile_X0E_Y0B_lo_out[6],Tile_X0E_Y0B_hi_out[6:5],Tile_X0E_Y0B_hi_out[5],Tile_X0E_Y0B_lo_out[4:3],Tile_X0E_Y0B_lo_out[3:2],Tile_X0E_Y0B_lo_out[2],Tile_X0E_Y0B_hi_out[2],Tile_X0E_Y0B_lo_out[1],Tile_X0E_Y0B_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X0E_Y0B_tile_id (
    .in(Tile_X0E_Y0B_tile_id_in),
    .out(Tile_X0E_Y0B_tile_id_out)
);
Tile_PE Tile_X0E_Y0C (
    .SB_T0_EAST_SB_IN_B1(Tile_X0F_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0F_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0E_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0E_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0E_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0E_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0E_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0E_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0E_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0E_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0E_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0E_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0D_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0D_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0E_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0E_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0F_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0F_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0E_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0E_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0E_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0E_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0E_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0E_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0E_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0E_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0E_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0E_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0D_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0D_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0E_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0E_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0F_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0F_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0E_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0E_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0E_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0E_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0E_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0E_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0E_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0E_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0E_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0E_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0D_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0D_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0E_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0E_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0F_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0F_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0E_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0E_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0E_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0E_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0E_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0E_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0E_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0E_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0E_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0E_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0D_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0D_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0E_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0E_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0F_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0F_Y0C_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0E_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0E_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0E_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0E_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0E_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0E_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0E_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0E_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0E_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0E_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0D_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0D_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0E_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0E_Y0C_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y0B_clk_out),
    .clk_out(Tile_X0E_Y0C_clk_out),
    .clk_pass_through(Tile_X0E_Y0B_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0E_Y0C_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0E_Y0C_clk_pass_through_out_right),
    .config_config_addr(Tile_X0E_Y0B_config_out_config_addr),
    .config_config_data(Tile_X0E_Y0B_config_out_config_data),
    .config_out_config_addr(Tile_X0E_Y0C_config_out_config_addr),
    .config_out_config_data(Tile_X0E_Y0C_config_out_config_data),
    .config_out_read(Tile_X0E_Y0C_config_out_read),
    .config_out_write(Tile_X0E_Y0C_config_out_write),
    .config_read(Tile_X0E_Y0B_config_out_read),
    .config_write(Tile_X0E_Y0B_config_out_write),
    .hi(Tile_X0E_Y0C_hi_unq1),
    .lo(Tile_X0E_Y0C_lo_unq1),
    .read_config_data(Tile_X0E_Y0C_read_config_data),
    .read_config_data_in(Tile_X0E_Y0B_read_config_data),
    .reset(Tile_X0E_Y0B_reset_out),
    .reset_out(Tile_X0E_Y0C_reset_out),
    .stall(Tile_X0E_Y0B_stall_out),
    .stall_out(Tile_X0E_Y0C_stall_out),
    .tile_id(Tile_X0E_Y0C_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0E_Y0C_hi (
    .in(Tile_X0E_Y0C_hi_unq1),
    .out(Tile_X0E_Y0C_hi_out)
);
mantle_wire__typeBit8 Tile_X0E_Y0C_lo (
    .in(Tile_X0E_Y0C_lo_unq1),
    .out(Tile_X0E_Y0C_lo_out)
);
wire [15:0] Tile_X0E_Y0C_tile_id_out;
assign Tile_X0E_Y0C_tile_id_out = {Tile_X0E_Y0C_lo_out[7],Tile_X0E_Y0C_lo_out[7:6],Tile_X0E_Y0C_lo_out[6],Tile_X0E_Y0C_hi_out[6:5],Tile_X0E_Y0C_hi_out[5],Tile_X0E_Y0C_lo_out[4:3],Tile_X0E_Y0C_lo_out[3:2],Tile_X0E_Y0C_lo_out[2],Tile_X0E_Y0C_hi_out[2:1],Tile_X0E_Y0C_lo_out[0],Tile_X0E_Y0C_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0E_Y0C_tile_id (
    .in(Tile_X0E_Y0C_tile_id_in),
    .out(Tile_X0E_Y0C_tile_id_out)
);
Tile_PE Tile_X0E_Y0D (
    .SB_T0_EAST_SB_IN_B1(Tile_X0F_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0F_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0E_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0E_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0E_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0E_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0E_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0E_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0E_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0E_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0E_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0E_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0D_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0D_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0E_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0E_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0F_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0F_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0E_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0E_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0E_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0E_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0E_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0E_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0E_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0E_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0E_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0E_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0D_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0D_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0E_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0E_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0F_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0F_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0E_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0E_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0E_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0E_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0E_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0E_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0E_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0E_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0E_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0E_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0D_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0D_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0E_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0E_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0F_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0F_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0E_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0E_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0E_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0E_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0E_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0E_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0E_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0E_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0E_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0E_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0D_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0D_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0E_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0E_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0F_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0F_Y0D_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0E_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0E_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0E_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0E_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0E_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0E_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0E_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0E_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0E_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0E_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0D_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0D_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0E_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0E_Y0D_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y0C_clk_out),
    .clk_out(Tile_X0E_Y0D_clk_out),
    .clk_pass_through(Tile_X0E_Y0C_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0E_Y0D_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0E_Y0D_clk_pass_through_out_right),
    .config_config_addr(Tile_X0E_Y0C_config_out_config_addr),
    .config_config_data(Tile_X0E_Y0C_config_out_config_data),
    .config_out_config_addr(Tile_X0E_Y0D_config_out_config_addr),
    .config_out_config_data(Tile_X0E_Y0D_config_out_config_data),
    .config_out_read(Tile_X0E_Y0D_config_out_read),
    .config_out_write(Tile_X0E_Y0D_config_out_write),
    .config_read(Tile_X0E_Y0C_config_out_read),
    .config_write(Tile_X0E_Y0C_config_out_write),
    .hi(Tile_X0E_Y0D_hi_unq1),
    .lo(Tile_X0E_Y0D_lo_unq1),
    .read_config_data(Tile_X0E_Y0D_read_config_data),
    .read_config_data_in(Tile_X0E_Y0C_read_config_data),
    .reset(Tile_X0E_Y0C_reset_out),
    .reset_out(Tile_X0E_Y0D_reset_out),
    .stall(Tile_X0E_Y0C_stall_out),
    .stall_out(Tile_X0E_Y0D_stall_out),
    .tile_id(Tile_X0E_Y0D_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0E_Y0D_hi (
    .in(Tile_X0E_Y0D_hi_unq1),
    .out(Tile_X0E_Y0D_hi_out)
);
mantle_wire__typeBit8 Tile_X0E_Y0D_lo (
    .in(Tile_X0E_Y0D_lo_unq1),
    .out(Tile_X0E_Y0D_lo_out)
);
wire [15:0] Tile_X0E_Y0D_tile_id_out;
assign Tile_X0E_Y0D_tile_id_out = {Tile_X0E_Y0D_lo_out[7],Tile_X0E_Y0D_lo_out[7:6],Tile_X0E_Y0D_lo_out[6],Tile_X0E_Y0D_hi_out[6:5],Tile_X0E_Y0D_hi_out[5],Tile_X0E_Y0D_lo_out[4:3],Tile_X0E_Y0D_lo_out[3:2],Tile_X0E_Y0D_lo_out[2],Tile_X0E_Y0D_hi_out[2:1],Tile_X0E_Y0D_lo_out[0],Tile_X0E_Y0D_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X0E_Y0D_tile_id (
    .in(Tile_X0E_Y0D_tile_id_in),
    .out(Tile_X0E_Y0D_tile_id_out)
);
Tile_PE Tile_X0E_Y0E (
    .SB_T0_EAST_SB_IN_B1(Tile_X0F_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0F_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0E_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0E_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0E_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0E_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0E_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0E_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0E_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0E_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0E_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0E_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0D_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0D_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0E_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0E_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0F_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0F_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0E_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0E_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0E_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0E_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0E_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0E_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0E_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0E_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0E_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0E_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0D_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0D_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0E_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0E_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0F_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0F_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0E_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0E_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0E_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0E_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0E_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0E_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0E_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0E_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0E_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0E_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0D_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0D_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0E_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0E_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0F_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0F_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0E_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0E_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0E_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0E_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0E_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0E_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0E_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0E_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0E_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0E_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0D_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0D_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0E_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0E_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0F_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0F_Y0E_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0E_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0E_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0E_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0E_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0E_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0E_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0E_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0E_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0E_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0E_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0D_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0D_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0E_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0E_Y0E_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y0D_clk_out),
    .clk_out(Tile_X0E_Y0E_clk_out),
    .clk_pass_through(Tile_X0E_Y0D_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0E_Y0E_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0E_Y0E_clk_pass_through_out_right),
    .config_config_addr(Tile_X0E_Y0D_config_out_config_addr),
    .config_config_data(Tile_X0E_Y0D_config_out_config_data),
    .config_out_config_addr(Tile_X0E_Y0E_config_out_config_addr),
    .config_out_config_data(Tile_X0E_Y0E_config_out_config_data),
    .config_out_read(Tile_X0E_Y0E_config_out_read),
    .config_out_write(Tile_X0E_Y0E_config_out_write),
    .config_read(Tile_X0E_Y0D_config_out_read),
    .config_write(Tile_X0E_Y0D_config_out_write),
    .hi(Tile_X0E_Y0E_hi_unq1),
    .lo(Tile_X0E_Y0E_lo_unq1),
    .read_config_data(Tile_X0E_Y0E_read_config_data),
    .read_config_data_in(Tile_X0E_Y0D_read_config_data),
    .reset(Tile_X0E_Y0D_reset_out),
    .reset_out(Tile_X0E_Y0E_reset_out),
    .stall(Tile_X0E_Y0D_stall_out),
    .stall_out(Tile_X0E_Y0E_stall_out),
    .tile_id(Tile_X0E_Y0E_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0E_Y0E_hi (
    .in(Tile_X0E_Y0E_hi_unq1),
    .out(Tile_X0E_Y0E_hi_out)
);
mantle_wire__typeBit8 Tile_X0E_Y0E_lo (
    .in(Tile_X0E_Y0E_lo_unq1),
    .out(Tile_X0E_Y0E_lo_out)
);
wire [15:0] Tile_X0E_Y0E_tile_id_out;
assign Tile_X0E_Y0E_tile_id_out = {Tile_X0E_Y0E_lo_out[7],Tile_X0E_Y0E_lo_out[7:6],Tile_X0E_Y0E_lo_out[6],Tile_X0E_Y0E_hi_out[6:5],Tile_X0E_Y0E_hi_out[5],Tile_X0E_Y0E_lo_out[4:3],Tile_X0E_Y0E_lo_out[3:2],Tile_X0E_Y0E_lo_out[2],Tile_X0E_Y0E_hi_out[2:1],Tile_X0E_Y0E_hi_out[1],Tile_X0E_Y0E_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0E_Y0E_tile_id (
    .in(Tile_X0E_Y0E_tile_id_in),
    .out(Tile_X0E_Y0E_tile_id_out)
);
Tile_PE Tile_X0E_Y0F (
    .SB_T0_EAST_SB_IN_B1(Tile_X0F_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0F_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0E_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0E_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0E_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0E_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0E_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0E_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0E_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0E_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0E_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0E_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0D_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0D_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0E_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0E_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0F_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0F_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0E_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0E_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0E_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0E_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0E_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0E_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0E_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0E_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0E_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0E_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0D_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0D_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0E_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0E_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0F_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0F_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0E_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0E_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0E_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0E_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0E_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0E_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0E_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0E_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0E_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0E_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0D_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0D_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0E_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0E_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0F_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0F_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0E_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0E_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0E_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0E_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0E_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0E_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0E_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0E_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0E_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0E_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0D_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0D_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0E_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0E_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0F_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0F_Y0F_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0E_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0E_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0E_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0E_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0E_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0E_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0E_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0E_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0E_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0E_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0D_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0D_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0E_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0E_Y0F_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y0E_clk_out),
    .clk_out(Tile_X0E_Y0F_clk_out),
    .clk_pass_through(Tile_X0E_Y0E_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0E_Y0F_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0E_Y0F_clk_pass_through_out_right),
    .config_config_addr(Tile_X0E_Y0E_config_out_config_addr),
    .config_config_data(Tile_X0E_Y0E_config_out_config_data),
    .config_out_config_addr(Tile_X0E_Y0F_config_out_config_addr),
    .config_out_config_data(Tile_X0E_Y0F_config_out_config_data),
    .config_out_read(Tile_X0E_Y0F_config_out_read),
    .config_out_write(Tile_X0E_Y0F_config_out_write),
    .config_read(Tile_X0E_Y0E_config_out_read),
    .config_write(Tile_X0E_Y0E_config_out_write),
    .hi(Tile_X0E_Y0F_hi_unq1),
    .lo(Tile_X0E_Y0F_lo_unq1),
    .read_config_data(Tile_X0E_Y0F_read_config_data),
    .read_config_data_in(Tile_X0E_Y0E_read_config_data),
    .reset(Tile_X0E_Y0E_reset_out),
    .reset_out(Tile_X0E_Y0F_reset_out),
    .stall(Tile_X0E_Y0E_stall_out),
    .stall_out(Tile_X0E_Y0F_stall_out),
    .tile_id(Tile_X0E_Y0F_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0E_Y0F_hi (
    .in(Tile_X0E_Y0F_hi_unq1),
    .out(Tile_X0E_Y0F_hi_out)
);
mantle_wire__typeBit8 Tile_X0E_Y0F_lo (
    .in(Tile_X0E_Y0F_lo_unq1),
    .out(Tile_X0E_Y0F_lo_out)
);
wire [15:0] Tile_X0E_Y0F_tile_id_out;
assign Tile_X0E_Y0F_tile_id_out = {Tile_X0E_Y0F_lo_out[7],Tile_X0E_Y0F_lo_out[7:6],Tile_X0E_Y0F_lo_out[6],Tile_X0E_Y0F_hi_out[6:5],Tile_X0E_Y0F_hi_out[5],Tile_X0E_Y0F_lo_out[4:3],Tile_X0E_Y0F_lo_out[3:2],Tile_X0E_Y0F_lo_out[2],Tile_X0E_Y0F_hi_out[2:1],Tile_X0E_Y0F_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X0E_Y0F_tile_id (
    .in(Tile_X0E_Y0F_tile_id_in),
    .out(Tile_X0E_Y0F_tile_id_out)
);
Tile_PE Tile_X0E_Y10 (
    .SB_T0_EAST_SB_IN_B1(Tile_X0F_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_EAST_SB_IN_B16(Tile_X0F_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0E_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0E_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0E_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0E_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0E_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0E_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T0_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0E_Y10_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0E_Y10_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0D_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0D_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0E_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0E_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(Tile_X0F_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_EAST_SB_IN_B16(Tile_X0F_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0E_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0E_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0E_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0E_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0E_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0E_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T1_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0E_Y10_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0E_Y10_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0D_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0D_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0E_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0E_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(Tile_X0F_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_EAST_SB_IN_B16(Tile_X0F_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0E_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0E_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0E_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0E_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0E_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0E_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T2_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0E_Y10_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0E_Y10_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0D_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0D_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0E_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0E_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(Tile_X0F_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_EAST_SB_IN_B16(Tile_X0F_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0E_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0E_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0E_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0E_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0E_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0E_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T3_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0E_Y10_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0E_Y10_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0D_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0D_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0E_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0E_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(Tile_X0F_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_EAST_SB_IN_B16(Tile_X0F_Y10_SB_T4_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0E_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0E_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0E_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0E_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0E_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0E_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T4_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0E_Y10_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0E_Y10_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0D_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0D_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0E_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0E_Y10_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y0F_clk_out),
    .clk_out(Tile_X0E_Y10_clk_out),
    .clk_pass_through(Tile_X0E_Y0F_clk_pass_through_out_bot),
    .clk_pass_through_out_bot(Tile_X0E_Y10_clk_pass_through_out_bot),
    .clk_pass_through_out_right(Tile_X0E_Y10_clk_pass_through_out_right),
    .config_config_addr(Tile_X0E_Y0F_config_out_config_addr),
    .config_config_data(Tile_X0E_Y0F_config_out_config_data),
    .config_out_config_addr(Tile_X0E_Y10_config_out_config_addr),
    .config_out_config_data(Tile_X0E_Y10_config_out_config_data),
    .config_out_read(Tile_X0E_Y10_config_out_read),
    .config_out_write(Tile_X0E_Y10_config_out_write),
    .config_read(Tile_X0E_Y0F_config_out_read),
    .config_write(Tile_X0E_Y0F_config_out_write),
    .hi(Tile_X0E_Y10_hi_unq1),
    .lo(Tile_X0E_Y10_lo_unq1),
    .read_config_data(Tile_X0E_Y10_read_config_data),
    .read_config_data_in(Tile_X0E_Y0F_read_config_data),
    .reset(Tile_X0E_Y0F_reset_out),
    .reset_out(Tile_X0E_Y10_reset_out),
    .stall(Tile_X0E_Y0F_stall_out),
    .stall_out(Tile_X0E_Y10_stall_out),
    .tile_id(Tile_X0E_Y10_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0E_Y10_hi (
    .in(Tile_X0E_Y10_hi_unq1),
    .out(Tile_X0E_Y10_hi_out)
);
mantle_wire__typeBit8 Tile_X0E_Y10_lo (
    .in(Tile_X0E_Y10_lo_unq1),
    .out(Tile_X0E_Y10_lo_out)
);
wire [15:0] Tile_X0E_Y10_tile_id_out;
assign Tile_X0E_Y10_tile_id_out = {Tile_X0E_Y10_lo_out[7],Tile_X0E_Y10_lo_out[7:6],Tile_X0E_Y10_lo_out[6],Tile_X0E_Y10_hi_out[6:5],Tile_X0E_Y10_hi_out[5],Tile_X0E_Y10_lo_out[4:3],Tile_X0E_Y10_lo_out[3:2],Tile_X0E_Y10_hi_out[2],Tile_X0E_Y10_lo_out[1],Tile_X0E_Y10_lo_out[1:0],Tile_X0E_Y10_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0E_Y10_tile_id (
    .in(Tile_X0E_Y10_tile_id_in),
    .out(Tile_X0E_Y10_tile_id_out)
);
wire [15:0] Tile_X0F_Y00_tile_id;
assign Tile_X0F_Y00_tile_id = {Tile_X0F_Y00_lo[7],Tile_X0F_Y00_lo[7:6],Tile_X0F_Y00_lo[6],Tile_X0F_Y00_hi[6:5],Tile_X0F_Y00_hi[5:4],Tile_X0F_Y00_lo[3],Tile_X0F_Y00_lo[3:2],Tile_X0F_Y00_lo[2:1],Tile_X0F_Y00_lo[1:0],Tile_X0F_Y00_lo[0]};
Tile_io_core Tile_X0F_Y00 (
    .tile_id(Tile_X0F_Y00_tile_id),
    .glb2io_1(glb2io_1_X0F_Y00),
    .f2io_1(Tile_X0F_Y01_SB_T0_NORTH_SB_OUT_B1),
    .io2glb_1(Tile_X0F_Y00_io2glb_1),
    .io2f_1(Tile_X0F_Y00_io2f_1),
    .glb2io_16(glb2io_16_X0F_Y00),
    .f2io_16(Tile_X0F_Y01_SB_T0_NORTH_SB_OUT_B16),
    .io2glb_16(Tile_X0F_Y00_io2glb_16),
    .io2f_16(Tile_X0F_Y00_io2f_16),
    .hi(Tile_X0F_Y00_hi),
    .lo(Tile_X0F_Y00_lo)
);
Tile_MemCore Tile_X0F_Y01 (
    .SB_T0_EAST_SB_IN_B1(const_0_1_out),
    .SB_T0_EAST_SB_IN_B16(const_0_16_out),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0F_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0F_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0F_Y00_io2f_1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0F_Y00_io2f_16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0F_Y01_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0F_Y01_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0F_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0F_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0F_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0F_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0E_Y01_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0E_Y01_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0F_Y01_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0F_Y01_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(const_0_1_out),
    .SB_T1_EAST_SB_IN_B16(const_0_16_out),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0F_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0F_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0F_Y00_io2f_1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0F_Y00_io2f_16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0F_Y01_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0F_Y01_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0F_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0F_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0F_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0F_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0E_Y01_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0E_Y01_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0F_Y01_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0F_Y01_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(const_0_1_out),
    .SB_T2_EAST_SB_IN_B16(const_0_16_out),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0F_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0F_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0F_Y00_io2f_1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0F_Y00_io2f_16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0F_Y01_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0F_Y01_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0F_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0F_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0F_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0F_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0E_Y01_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0E_Y01_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0F_Y01_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0F_Y01_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(const_0_1_out),
    .SB_T3_EAST_SB_IN_B16(const_0_16_out),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0F_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0F_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0F_Y00_io2f_1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0F_Y00_io2f_16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0F_Y01_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0F_Y01_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0F_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0F_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0F_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0F_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0E_Y01_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0E_Y01_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0F_Y01_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0F_Y01_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(const_0_1_out),
    .SB_T4_EAST_SB_IN_B16(const_0_16_out),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0F_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0F_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0F_Y00_io2f_1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0F_Y00_io2f_16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0F_Y01_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0F_Y01_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0F_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0F_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0F_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0F_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0E_Y01_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0E_Y01_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0F_Y01_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0F_Y01_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y01_clk_pass_through_out_right),
    .clk_out(Tile_X0F_Y01_clk_out),
    .config_config_addr(config_15_config_addr),
    .config_config_data(config_15_config_data),
    .config_out_config_addr(Tile_X0F_Y01_config_out_config_addr),
    .config_out_config_data(Tile_X0F_Y01_config_out_config_data),
    .config_out_read(Tile_X0F_Y01_config_out_read),
    .config_out_write(Tile_X0F_Y01_config_out_write),
    .config_read(config_15_read),
    .config_write(config_15_write),
    .hi(Tile_X0F_Y01_hi_unq1),
    .lo(Tile_X0F_Y01_lo_unq1),
    .read_config_data(Tile_X0F_Y01_read_config_data),
    .read_config_data_in(const_0_32_out),
    .reset(reset),
    .reset_out(Tile_X0F_Y01_reset_out),
    .stall(stall[15]),
    .stall_out(Tile_X0F_Y01_stall_out),
    .tile_id(Tile_X0F_Y01_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0F_Y01_hi (
    .in(Tile_X0F_Y01_hi_unq1),
    .out(Tile_X0F_Y01_hi_out)
);
mantle_wire__typeBit8 Tile_X0F_Y01_lo (
    .in(Tile_X0F_Y01_lo_unq1),
    .out(Tile_X0F_Y01_lo_out)
);
wire [15:0] Tile_X0F_Y01_tile_id_out;
assign Tile_X0F_Y01_tile_id_out = {Tile_X0F_Y01_lo_out[7],Tile_X0F_Y01_lo_out[7:6],Tile_X0F_Y01_lo_out[6],Tile_X0F_Y01_hi_out[6:5],Tile_X0F_Y01_hi_out[5:4],Tile_X0F_Y01_lo_out[3],Tile_X0F_Y01_lo_out[3:2],Tile_X0F_Y01_lo_out[2:1],Tile_X0F_Y01_lo_out[1:0],Tile_X0F_Y01_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X0F_Y01_tile_id (
    .in(Tile_X0F_Y01_tile_id_in),
    .out(Tile_X0F_Y01_tile_id_out)
);
Tile_MemCore Tile_X0F_Y02 (
    .SB_T0_EAST_SB_IN_B1(const_0_1_out),
    .SB_T0_EAST_SB_IN_B16(const_0_16_out),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0F_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0F_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0F_Y01_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0F_Y01_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0F_Y02_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0F_Y02_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0F_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0F_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0F_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0F_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0E_Y02_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0E_Y02_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0F_Y02_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0F_Y02_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(const_0_1_out),
    .SB_T1_EAST_SB_IN_B16(const_0_16_out),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0F_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0F_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0F_Y01_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0F_Y01_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0F_Y02_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0F_Y02_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0F_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0F_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0F_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0F_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0E_Y02_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0E_Y02_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0F_Y02_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0F_Y02_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(const_0_1_out),
    .SB_T2_EAST_SB_IN_B16(const_0_16_out),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0F_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0F_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0F_Y01_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0F_Y01_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0F_Y02_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0F_Y02_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0F_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0F_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0F_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0F_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0E_Y02_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0E_Y02_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0F_Y02_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0F_Y02_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(const_0_1_out),
    .SB_T3_EAST_SB_IN_B16(const_0_16_out),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0F_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0F_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0F_Y01_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0F_Y01_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0F_Y02_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0F_Y02_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0F_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0F_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0F_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0F_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0E_Y02_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0E_Y02_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0F_Y02_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0F_Y02_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(const_0_1_out),
    .SB_T4_EAST_SB_IN_B16(const_0_16_out),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0F_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0F_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0F_Y01_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0F_Y01_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0F_Y02_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0F_Y02_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0F_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0F_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0F_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0F_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0E_Y02_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0E_Y02_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0F_Y02_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0F_Y02_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y02_clk_pass_through_out_right),
    .clk_out(Tile_X0F_Y02_clk_out),
    .config_config_addr(Tile_X0F_Y01_config_out_config_addr),
    .config_config_data(Tile_X0F_Y01_config_out_config_data),
    .config_out_config_addr(Tile_X0F_Y02_config_out_config_addr),
    .config_out_config_data(Tile_X0F_Y02_config_out_config_data),
    .config_out_read(Tile_X0F_Y02_config_out_read),
    .config_out_write(Tile_X0F_Y02_config_out_write),
    .config_read(Tile_X0F_Y01_config_out_read),
    .config_write(Tile_X0F_Y01_config_out_write),
    .hi(Tile_X0F_Y02_hi_unq1),
    .lo(Tile_X0F_Y02_lo_unq1),
    .read_config_data(Tile_X0F_Y02_read_config_data),
    .read_config_data_in(Tile_X0F_Y01_read_config_data),
    .reset(Tile_X0F_Y01_reset_out),
    .reset_out(Tile_X0F_Y02_reset_out),
    .stall(Tile_X0F_Y01_stall_out),
    .stall_out(Tile_X0F_Y02_stall_out),
    .tile_id(Tile_X0F_Y02_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0F_Y02_hi (
    .in(Tile_X0F_Y02_hi_unq1),
    .out(Tile_X0F_Y02_hi_out)
);
mantle_wire__typeBit8 Tile_X0F_Y02_lo (
    .in(Tile_X0F_Y02_lo_unq1),
    .out(Tile_X0F_Y02_lo_out)
);
wire [15:0] Tile_X0F_Y02_tile_id_out;
assign Tile_X0F_Y02_tile_id_out = {Tile_X0F_Y02_lo_out[7],Tile_X0F_Y02_lo_out[7:6],Tile_X0F_Y02_lo_out[6],Tile_X0F_Y02_hi_out[6:5],Tile_X0F_Y02_hi_out[5:4],Tile_X0F_Y02_lo_out[3],Tile_X0F_Y02_lo_out[3:2],Tile_X0F_Y02_lo_out[2:1],Tile_X0F_Y02_lo_out[1],Tile_X0F_Y02_hi_out[1],Tile_X0F_Y02_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0F_Y02_tile_id (
    .in(Tile_X0F_Y02_tile_id_in),
    .out(Tile_X0F_Y02_tile_id_out)
);
Tile_MemCore Tile_X0F_Y03 (
    .SB_T0_EAST_SB_IN_B1(const_0_1_out),
    .SB_T0_EAST_SB_IN_B16(const_0_16_out),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0F_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0F_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0F_Y02_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0F_Y02_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0F_Y03_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0F_Y03_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0F_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0F_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0F_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0F_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0E_Y03_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0E_Y03_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0F_Y03_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0F_Y03_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(const_0_1_out),
    .SB_T1_EAST_SB_IN_B16(const_0_16_out),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0F_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0F_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0F_Y02_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0F_Y02_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0F_Y03_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0F_Y03_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0F_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0F_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0F_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0F_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0E_Y03_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0E_Y03_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0F_Y03_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0F_Y03_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(const_0_1_out),
    .SB_T2_EAST_SB_IN_B16(const_0_16_out),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0F_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0F_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0F_Y02_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0F_Y02_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0F_Y03_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0F_Y03_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0F_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0F_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0F_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0F_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0E_Y03_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0E_Y03_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0F_Y03_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0F_Y03_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(const_0_1_out),
    .SB_T3_EAST_SB_IN_B16(const_0_16_out),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0F_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0F_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0F_Y02_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0F_Y02_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0F_Y03_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0F_Y03_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0F_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0F_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0F_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0F_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0E_Y03_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0E_Y03_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0F_Y03_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0F_Y03_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(const_0_1_out),
    .SB_T4_EAST_SB_IN_B16(const_0_16_out),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0F_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0F_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0F_Y02_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0F_Y02_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0F_Y03_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0F_Y03_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0F_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0F_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0F_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0F_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0E_Y03_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0E_Y03_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0F_Y03_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0F_Y03_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y03_clk_pass_through_out_right),
    .clk_out(Tile_X0F_Y03_clk_out),
    .config_config_addr(Tile_X0F_Y02_config_out_config_addr),
    .config_config_data(Tile_X0F_Y02_config_out_config_data),
    .config_out_config_addr(Tile_X0F_Y03_config_out_config_addr),
    .config_out_config_data(Tile_X0F_Y03_config_out_config_data),
    .config_out_read(Tile_X0F_Y03_config_out_read),
    .config_out_write(Tile_X0F_Y03_config_out_write),
    .config_read(Tile_X0F_Y02_config_out_read),
    .config_write(Tile_X0F_Y02_config_out_write),
    .hi(Tile_X0F_Y03_hi_unq1),
    .lo(Tile_X0F_Y03_lo_unq1),
    .read_config_data(Tile_X0F_Y03_read_config_data),
    .read_config_data_in(Tile_X0F_Y02_read_config_data),
    .reset(Tile_X0F_Y02_reset_out),
    .reset_out(Tile_X0F_Y03_reset_out),
    .stall(Tile_X0F_Y02_stall_out),
    .stall_out(Tile_X0F_Y03_stall_out),
    .tile_id(Tile_X0F_Y03_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0F_Y03_hi (
    .in(Tile_X0F_Y03_hi_unq1),
    .out(Tile_X0F_Y03_hi_out)
);
mantle_wire__typeBit8 Tile_X0F_Y03_lo (
    .in(Tile_X0F_Y03_lo_unq1),
    .out(Tile_X0F_Y03_lo_out)
);
wire [15:0] Tile_X0F_Y03_tile_id_out;
assign Tile_X0F_Y03_tile_id_out = {Tile_X0F_Y03_lo_out[7],Tile_X0F_Y03_lo_out[7:6],Tile_X0F_Y03_lo_out[6],Tile_X0F_Y03_hi_out[6:5],Tile_X0F_Y03_hi_out[5:4],Tile_X0F_Y03_lo_out[3],Tile_X0F_Y03_lo_out[3:2],Tile_X0F_Y03_lo_out[2:1],Tile_X0F_Y03_lo_out[1],Tile_X0F_Y03_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X0F_Y03_tile_id (
    .in(Tile_X0F_Y03_tile_id_in),
    .out(Tile_X0F_Y03_tile_id_out)
);
Tile_MemCore Tile_X0F_Y04 (
    .SB_T0_EAST_SB_IN_B1(const_0_1_out),
    .SB_T0_EAST_SB_IN_B16(const_0_16_out),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0F_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0F_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0F_Y03_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0F_Y03_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0F_Y04_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0F_Y04_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0F_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0F_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0F_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0F_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0E_Y04_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0E_Y04_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0F_Y04_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0F_Y04_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(const_0_1_out),
    .SB_T1_EAST_SB_IN_B16(const_0_16_out),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0F_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0F_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0F_Y03_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0F_Y03_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0F_Y04_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0F_Y04_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0F_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0F_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0F_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0F_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0E_Y04_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0E_Y04_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0F_Y04_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0F_Y04_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(const_0_1_out),
    .SB_T2_EAST_SB_IN_B16(const_0_16_out),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0F_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0F_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0F_Y03_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0F_Y03_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0F_Y04_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0F_Y04_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0F_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0F_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0F_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0F_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0E_Y04_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0E_Y04_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0F_Y04_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0F_Y04_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(const_0_1_out),
    .SB_T3_EAST_SB_IN_B16(const_0_16_out),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0F_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0F_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0F_Y03_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0F_Y03_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0F_Y04_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0F_Y04_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0F_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0F_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0F_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0F_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0E_Y04_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0E_Y04_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0F_Y04_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0F_Y04_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(const_0_1_out),
    .SB_T4_EAST_SB_IN_B16(const_0_16_out),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0F_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0F_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0F_Y03_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0F_Y03_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0F_Y04_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0F_Y04_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0F_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0F_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0F_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0F_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0E_Y04_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0E_Y04_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0F_Y04_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0F_Y04_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y04_clk_pass_through_out_right),
    .clk_out(Tile_X0F_Y04_clk_out),
    .config_config_addr(Tile_X0F_Y03_config_out_config_addr),
    .config_config_data(Tile_X0F_Y03_config_out_config_data),
    .config_out_config_addr(Tile_X0F_Y04_config_out_config_addr),
    .config_out_config_data(Tile_X0F_Y04_config_out_config_data),
    .config_out_read(Tile_X0F_Y04_config_out_read),
    .config_out_write(Tile_X0F_Y04_config_out_write),
    .config_read(Tile_X0F_Y03_config_out_read),
    .config_write(Tile_X0F_Y03_config_out_write),
    .hi(Tile_X0F_Y04_hi_unq1),
    .lo(Tile_X0F_Y04_lo_unq1),
    .read_config_data(Tile_X0F_Y04_read_config_data),
    .read_config_data_in(Tile_X0F_Y03_read_config_data),
    .reset(Tile_X0F_Y03_reset_out),
    .reset_out(Tile_X0F_Y04_reset_out),
    .stall(Tile_X0F_Y03_stall_out),
    .stall_out(Tile_X0F_Y04_stall_out),
    .tile_id(Tile_X0F_Y04_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0F_Y04_hi (
    .in(Tile_X0F_Y04_hi_unq1),
    .out(Tile_X0F_Y04_hi_out)
);
mantle_wire__typeBit8 Tile_X0F_Y04_lo (
    .in(Tile_X0F_Y04_lo_unq1),
    .out(Tile_X0F_Y04_lo_out)
);
wire [15:0] Tile_X0F_Y04_tile_id_out;
assign Tile_X0F_Y04_tile_id_out = {Tile_X0F_Y04_lo_out[7],Tile_X0F_Y04_lo_out[7:6],Tile_X0F_Y04_lo_out[6],Tile_X0F_Y04_hi_out[6:5],Tile_X0F_Y04_hi_out[5:4],Tile_X0F_Y04_lo_out[3],Tile_X0F_Y04_lo_out[3:2],Tile_X0F_Y04_lo_out[2:1],Tile_X0F_Y04_hi_out[1],Tile_X0F_Y04_lo_out[0],Tile_X0F_Y04_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0F_Y04_tile_id (
    .in(Tile_X0F_Y04_tile_id_in),
    .out(Tile_X0F_Y04_tile_id_out)
);
Tile_MemCore Tile_X0F_Y05 (
    .SB_T0_EAST_SB_IN_B1(const_0_1_out),
    .SB_T0_EAST_SB_IN_B16(const_0_16_out),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0F_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0F_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0F_Y04_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0F_Y04_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0F_Y05_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0F_Y05_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0F_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0F_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0F_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0F_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0E_Y05_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0E_Y05_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0F_Y05_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0F_Y05_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(const_0_1_out),
    .SB_T1_EAST_SB_IN_B16(const_0_16_out),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0F_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0F_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0F_Y04_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0F_Y04_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0F_Y05_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0F_Y05_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0F_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0F_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0F_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0F_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0E_Y05_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0E_Y05_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0F_Y05_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0F_Y05_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(const_0_1_out),
    .SB_T2_EAST_SB_IN_B16(const_0_16_out),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0F_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0F_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0F_Y04_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0F_Y04_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0F_Y05_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0F_Y05_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0F_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0F_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0F_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0F_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0E_Y05_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0E_Y05_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0F_Y05_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0F_Y05_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(const_0_1_out),
    .SB_T3_EAST_SB_IN_B16(const_0_16_out),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0F_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0F_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0F_Y04_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0F_Y04_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0F_Y05_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0F_Y05_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0F_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0F_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0F_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0F_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0E_Y05_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0E_Y05_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0F_Y05_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0F_Y05_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(const_0_1_out),
    .SB_T4_EAST_SB_IN_B16(const_0_16_out),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0F_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0F_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0F_Y04_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0F_Y04_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0F_Y05_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0F_Y05_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0F_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0F_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0F_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0F_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0E_Y05_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0E_Y05_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0F_Y05_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0F_Y05_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y05_clk_pass_through_out_right),
    .clk_out(Tile_X0F_Y05_clk_out),
    .config_config_addr(Tile_X0F_Y04_config_out_config_addr),
    .config_config_data(Tile_X0F_Y04_config_out_config_data),
    .config_out_config_addr(Tile_X0F_Y05_config_out_config_addr),
    .config_out_config_data(Tile_X0F_Y05_config_out_config_data),
    .config_out_read(Tile_X0F_Y05_config_out_read),
    .config_out_write(Tile_X0F_Y05_config_out_write),
    .config_read(Tile_X0F_Y04_config_out_read),
    .config_write(Tile_X0F_Y04_config_out_write),
    .hi(Tile_X0F_Y05_hi_unq1),
    .lo(Tile_X0F_Y05_lo_unq1),
    .read_config_data(Tile_X0F_Y05_read_config_data),
    .read_config_data_in(Tile_X0F_Y04_read_config_data),
    .reset(Tile_X0F_Y04_reset_out),
    .reset_out(Tile_X0F_Y05_reset_out),
    .stall(Tile_X0F_Y04_stall_out),
    .stall_out(Tile_X0F_Y05_stall_out),
    .tile_id(Tile_X0F_Y05_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0F_Y05_hi (
    .in(Tile_X0F_Y05_hi_unq1),
    .out(Tile_X0F_Y05_hi_out)
);
mantle_wire__typeBit8 Tile_X0F_Y05_lo (
    .in(Tile_X0F_Y05_lo_unq1),
    .out(Tile_X0F_Y05_lo_out)
);
wire [15:0] Tile_X0F_Y05_tile_id_out;
assign Tile_X0F_Y05_tile_id_out = {Tile_X0F_Y05_lo_out[7],Tile_X0F_Y05_lo_out[7:6],Tile_X0F_Y05_lo_out[6],Tile_X0F_Y05_hi_out[6:5],Tile_X0F_Y05_hi_out[5:4],Tile_X0F_Y05_lo_out[3],Tile_X0F_Y05_lo_out[3:2],Tile_X0F_Y05_lo_out[2:1],Tile_X0F_Y05_hi_out[1],Tile_X0F_Y05_lo_out[0],Tile_X0F_Y05_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X0F_Y05_tile_id (
    .in(Tile_X0F_Y05_tile_id_in),
    .out(Tile_X0F_Y05_tile_id_out)
);
Tile_MemCore Tile_X0F_Y06 (
    .SB_T0_EAST_SB_IN_B1(const_0_1_out),
    .SB_T0_EAST_SB_IN_B16(const_0_16_out),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0F_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0F_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0F_Y05_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0F_Y05_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0F_Y06_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0F_Y06_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0F_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0F_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0F_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0F_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0E_Y06_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0E_Y06_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0F_Y06_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0F_Y06_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(const_0_1_out),
    .SB_T1_EAST_SB_IN_B16(const_0_16_out),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0F_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0F_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0F_Y05_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0F_Y05_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0F_Y06_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0F_Y06_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0F_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0F_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0F_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0F_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0E_Y06_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0E_Y06_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0F_Y06_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0F_Y06_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(const_0_1_out),
    .SB_T2_EAST_SB_IN_B16(const_0_16_out),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0F_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0F_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0F_Y05_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0F_Y05_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0F_Y06_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0F_Y06_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0F_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0F_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0F_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0F_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0E_Y06_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0E_Y06_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0F_Y06_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0F_Y06_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(const_0_1_out),
    .SB_T3_EAST_SB_IN_B16(const_0_16_out),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0F_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0F_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0F_Y05_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0F_Y05_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0F_Y06_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0F_Y06_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0F_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0F_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0F_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0F_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0E_Y06_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0E_Y06_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0F_Y06_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0F_Y06_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(const_0_1_out),
    .SB_T4_EAST_SB_IN_B16(const_0_16_out),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0F_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0F_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0F_Y05_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0F_Y05_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0F_Y06_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0F_Y06_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0F_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0F_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0F_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0F_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0E_Y06_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0E_Y06_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0F_Y06_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0F_Y06_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y06_clk_pass_through_out_right),
    .clk_out(Tile_X0F_Y06_clk_out),
    .config_config_addr(Tile_X0F_Y05_config_out_config_addr),
    .config_config_data(Tile_X0F_Y05_config_out_config_data),
    .config_out_config_addr(Tile_X0F_Y06_config_out_config_addr),
    .config_out_config_data(Tile_X0F_Y06_config_out_config_data),
    .config_out_read(Tile_X0F_Y06_config_out_read),
    .config_out_write(Tile_X0F_Y06_config_out_write),
    .config_read(Tile_X0F_Y05_config_out_read),
    .config_write(Tile_X0F_Y05_config_out_write),
    .hi(Tile_X0F_Y06_hi_unq1),
    .lo(Tile_X0F_Y06_lo_unq1),
    .read_config_data(Tile_X0F_Y06_read_config_data),
    .read_config_data_in(Tile_X0F_Y05_read_config_data),
    .reset(Tile_X0F_Y05_reset_out),
    .reset_out(Tile_X0F_Y06_reset_out),
    .stall(Tile_X0F_Y05_stall_out),
    .stall_out(Tile_X0F_Y06_stall_out),
    .tile_id(Tile_X0F_Y06_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0F_Y06_hi (
    .in(Tile_X0F_Y06_hi_unq1),
    .out(Tile_X0F_Y06_hi_out)
);
mantle_wire__typeBit8 Tile_X0F_Y06_lo (
    .in(Tile_X0F_Y06_lo_unq1),
    .out(Tile_X0F_Y06_lo_out)
);
wire [15:0] Tile_X0F_Y06_tile_id_out;
assign Tile_X0F_Y06_tile_id_out = {Tile_X0F_Y06_lo_out[7],Tile_X0F_Y06_lo_out[7:6],Tile_X0F_Y06_lo_out[6],Tile_X0F_Y06_hi_out[6:5],Tile_X0F_Y06_hi_out[5:4],Tile_X0F_Y06_lo_out[3],Tile_X0F_Y06_lo_out[3:2],Tile_X0F_Y06_lo_out[2:1],Tile_X0F_Y06_hi_out[1],Tile_X0F_Y06_hi_out[1],Tile_X0F_Y06_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0F_Y06_tile_id (
    .in(Tile_X0F_Y06_tile_id_in),
    .out(Tile_X0F_Y06_tile_id_out)
);
Tile_MemCore Tile_X0F_Y07 (
    .SB_T0_EAST_SB_IN_B1(const_0_1_out),
    .SB_T0_EAST_SB_IN_B16(const_0_16_out),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0F_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0F_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0F_Y06_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0F_Y06_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0F_Y07_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0F_Y07_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0F_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0F_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0F_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0F_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0E_Y07_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0E_Y07_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0F_Y07_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0F_Y07_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(const_0_1_out),
    .SB_T1_EAST_SB_IN_B16(const_0_16_out),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0F_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0F_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0F_Y06_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0F_Y06_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0F_Y07_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0F_Y07_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0F_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0F_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0F_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0F_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0E_Y07_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0E_Y07_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0F_Y07_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0F_Y07_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(const_0_1_out),
    .SB_T2_EAST_SB_IN_B16(const_0_16_out),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0F_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0F_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0F_Y06_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0F_Y06_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0F_Y07_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0F_Y07_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0F_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0F_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0F_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0F_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0E_Y07_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0E_Y07_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0F_Y07_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0F_Y07_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(const_0_1_out),
    .SB_T3_EAST_SB_IN_B16(const_0_16_out),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0F_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0F_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0F_Y06_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0F_Y06_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0F_Y07_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0F_Y07_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0F_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0F_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0F_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0F_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0E_Y07_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0E_Y07_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0F_Y07_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0F_Y07_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(const_0_1_out),
    .SB_T4_EAST_SB_IN_B16(const_0_16_out),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0F_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0F_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0F_Y06_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0F_Y06_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0F_Y07_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0F_Y07_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0F_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0F_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0F_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0F_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0E_Y07_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0E_Y07_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0F_Y07_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0F_Y07_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y07_clk_pass_through_out_right),
    .clk_out(Tile_X0F_Y07_clk_out),
    .config_config_addr(Tile_X0F_Y06_config_out_config_addr),
    .config_config_data(Tile_X0F_Y06_config_out_config_data),
    .config_out_config_addr(Tile_X0F_Y07_config_out_config_addr),
    .config_out_config_data(Tile_X0F_Y07_config_out_config_data),
    .config_out_read(Tile_X0F_Y07_config_out_read),
    .config_out_write(Tile_X0F_Y07_config_out_write),
    .config_read(Tile_X0F_Y06_config_out_read),
    .config_write(Tile_X0F_Y06_config_out_write),
    .hi(Tile_X0F_Y07_hi_unq1),
    .lo(Tile_X0F_Y07_lo_unq1),
    .read_config_data(Tile_X0F_Y07_read_config_data),
    .read_config_data_in(Tile_X0F_Y06_read_config_data),
    .reset(Tile_X0F_Y06_reset_out),
    .reset_out(Tile_X0F_Y07_reset_out),
    .stall(Tile_X0F_Y06_stall_out),
    .stall_out(Tile_X0F_Y07_stall_out),
    .tile_id(Tile_X0F_Y07_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0F_Y07_hi (
    .in(Tile_X0F_Y07_hi_unq1),
    .out(Tile_X0F_Y07_hi_out)
);
mantle_wire__typeBit8 Tile_X0F_Y07_lo (
    .in(Tile_X0F_Y07_lo_unq1),
    .out(Tile_X0F_Y07_lo_out)
);
wire [15:0] Tile_X0F_Y07_tile_id_out;
assign Tile_X0F_Y07_tile_id_out = {Tile_X0F_Y07_lo_out[7],Tile_X0F_Y07_lo_out[7:6],Tile_X0F_Y07_lo_out[6],Tile_X0F_Y07_hi_out[6:5],Tile_X0F_Y07_hi_out[5:4],Tile_X0F_Y07_lo_out[3],Tile_X0F_Y07_lo_out[3:2],Tile_X0F_Y07_lo_out[2:1],Tile_X0F_Y07_hi_out[1],Tile_X0F_Y07_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X0F_Y07_tile_id (
    .in(Tile_X0F_Y07_tile_id_in),
    .out(Tile_X0F_Y07_tile_id_out)
);
Tile_MemCore Tile_X0F_Y08 (
    .SB_T0_EAST_SB_IN_B1(const_0_1_out),
    .SB_T0_EAST_SB_IN_B16(const_0_16_out),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0F_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0F_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0F_Y07_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0F_Y07_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0F_Y08_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0F_Y08_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0F_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0F_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0F_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0F_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0E_Y08_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0E_Y08_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0F_Y08_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0F_Y08_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(const_0_1_out),
    .SB_T1_EAST_SB_IN_B16(const_0_16_out),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0F_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0F_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0F_Y07_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0F_Y07_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0F_Y08_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0F_Y08_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0F_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0F_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0F_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0F_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0E_Y08_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0E_Y08_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0F_Y08_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0F_Y08_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(const_0_1_out),
    .SB_T2_EAST_SB_IN_B16(const_0_16_out),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0F_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0F_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0F_Y07_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0F_Y07_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0F_Y08_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0F_Y08_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0F_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0F_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0F_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0F_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0E_Y08_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0E_Y08_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0F_Y08_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0F_Y08_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(const_0_1_out),
    .SB_T3_EAST_SB_IN_B16(const_0_16_out),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0F_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0F_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0F_Y07_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0F_Y07_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0F_Y08_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0F_Y08_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0F_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0F_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0F_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0F_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0E_Y08_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0E_Y08_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0F_Y08_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0F_Y08_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(const_0_1_out),
    .SB_T4_EAST_SB_IN_B16(const_0_16_out),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0F_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0F_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0F_Y07_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0F_Y07_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0F_Y08_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0F_Y08_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0F_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0F_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0F_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0F_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0E_Y08_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0E_Y08_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0F_Y08_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0F_Y08_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y08_clk_pass_through_out_right),
    .clk_out(Tile_X0F_Y08_clk_out),
    .config_config_addr(Tile_X0F_Y07_config_out_config_addr),
    .config_config_data(Tile_X0F_Y07_config_out_config_data),
    .config_out_config_addr(Tile_X0F_Y08_config_out_config_addr),
    .config_out_config_data(Tile_X0F_Y08_config_out_config_data),
    .config_out_read(Tile_X0F_Y08_config_out_read),
    .config_out_write(Tile_X0F_Y08_config_out_write),
    .config_read(Tile_X0F_Y07_config_out_read),
    .config_write(Tile_X0F_Y07_config_out_write),
    .hi(Tile_X0F_Y08_hi_unq1),
    .lo(Tile_X0F_Y08_lo_unq1),
    .read_config_data(Tile_X0F_Y08_read_config_data),
    .read_config_data_in(Tile_X0F_Y07_read_config_data),
    .reset(Tile_X0F_Y07_reset_out),
    .reset_out(Tile_X0F_Y08_reset_out),
    .stall(Tile_X0F_Y07_stall_out),
    .stall_out(Tile_X0F_Y08_stall_out),
    .tile_id(Tile_X0F_Y08_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0F_Y08_hi (
    .in(Tile_X0F_Y08_hi_unq1),
    .out(Tile_X0F_Y08_hi_out)
);
mantle_wire__typeBit8 Tile_X0F_Y08_lo (
    .in(Tile_X0F_Y08_lo_unq1),
    .out(Tile_X0F_Y08_lo_out)
);
wire [15:0] Tile_X0F_Y08_tile_id_out;
assign Tile_X0F_Y08_tile_id_out = {Tile_X0F_Y08_lo_out[7],Tile_X0F_Y08_lo_out[7:6],Tile_X0F_Y08_lo_out[6],Tile_X0F_Y08_hi_out[6:5],Tile_X0F_Y08_hi_out[5:4],Tile_X0F_Y08_lo_out[3],Tile_X0F_Y08_lo_out[3:2],Tile_X0F_Y08_lo_out[2],Tile_X0F_Y08_hi_out[2],Tile_X0F_Y08_lo_out[1:0],Tile_X0F_Y08_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0F_Y08_tile_id (
    .in(Tile_X0F_Y08_tile_id_in),
    .out(Tile_X0F_Y08_tile_id_out)
);
Tile_MemCore Tile_X0F_Y09 (
    .SB_T0_EAST_SB_IN_B1(const_0_1_out),
    .SB_T0_EAST_SB_IN_B16(const_0_16_out),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0F_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0F_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0F_Y08_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0F_Y08_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0F_Y09_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0F_Y09_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0F_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0F_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0F_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0F_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0E_Y09_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0E_Y09_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0F_Y09_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0F_Y09_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(const_0_1_out),
    .SB_T1_EAST_SB_IN_B16(const_0_16_out),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0F_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0F_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0F_Y08_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0F_Y08_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0F_Y09_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0F_Y09_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0F_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0F_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0F_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0F_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0E_Y09_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0E_Y09_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0F_Y09_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0F_Y09_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(const_0_1_out),
    .SB_T2_EAST_SB_IN_B16(const_0_16_out),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0F_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0F_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0F_Y08_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0F_Y08_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0F_Y09_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0F_Y09_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0F_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0F_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0F_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0F_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0E_Y09_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0E_Y09_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0F_Y09_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0F_Y09_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(const_0_1_out),
    .SB_T3_EAST_SB_IN_B16(const_0_16_out),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0F_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0F_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0F_Y08_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0F_Y08_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0F_Y09_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0F_Y09_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0F_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0F_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0F_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0F_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0E_Y09_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0E_Y09_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0F_Y09_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0F_Y09_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(const_0_1_out),
    .SB_T4_EAST_SB_IN_B16(const_0_16_out),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0F_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0F_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0F_Y08_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0F_Y08_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0F_Y09_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0F_Y09_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0F_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0F_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0F_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0F_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0E_Y09_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0E_Y09_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0F_Y09_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0F_Y09_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y09_clk_pass_through_out_right),
    .clk_out(Tile_X0F_Y09_clk_out),
    .config_config_addr(ConfigPipeStage_inst15_config_out_config_addr),
    .config_config_data(ConfigPipeStage_inst15_config_out_config_data),
    .config_out_config_addr(Tile_X0F_Y09_config_out_config_addr),
    .config_out_config_data(Tile_X0F_Y09_config_out_config_data),
    .config_out_read(Tile_X0F_Y09_config_out_read),
    .config_out_write(Tile_X0F_Y09_config_out_write),
    .config_read(ConfigPipeStage_inst15_config_out_read),
    .config_write(ConfigPipeStage_inst15_config_out_write),
    .hi(Tile_X0F_Y09_hi_unq1),
    .lo(Tile_X0F_Y09_lo_unq1),
    .read_config_data(Tile_X0F_Y09_read_config_data),
    .read_config_data_in(Tile_X0F_Y08_read_config_data),
    .reset(Tile_X0F_Y08_reset_out),
    .reset_out(Tile_X0F_Y09_reset_out),
    .stall(Tile_X0F_Y08_stall_out),
    .stall_out(Tile_X0F_Y09_stall_out),
    .tile_id(Tile_X0F_Y09_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0F_Y09_hi (
    .in(Tile_X0F_Y09_hi_unq1),
    .out(Tile_X0F_Y09_hi_out)
);
mantle_wire__typeBit8 Tile_X0F_Y09_lo (
    .in(Tile_X0F_Y09_lo_unq1),
    .out(Tile_X0F_Y09_lo_out)
);
wire [15:0] Tile_X0F_Y09_tile_id_out;
assign Tile_X0F_Y09_tile_id_out = {Tile_X0F_Y09_lo_out[7],Tile_X0F_Y09_lo_out[7:6],Tile_X0F_Y09_lo_out[6],Tile_X0F_Y09_hi_out[6:5],Tile_X0F_Y09_hi_out[5:4],Tile_X0F_Y09_lo_out[3],Tile_X0F_Y09_lo_out[3:2],Tile_X0F_Y09_lo_out[2],Tile_X0F_Y09_hi_out[2],Tile_X0F_Y09_lo_out[1:0],Tile_X0F_Y09_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X0F_Y09_tile_id (
    .in(Tile_X0F_Y09_tile_id_in),
    .out(Tile_X0F_Y09_tile_id_out)
);
Tile_MemCore Tile_X0F_Y0A (
    .SB_T0_EAST_SB_IN_B1(const_0_1_out),
    .SB_T0_EAST_SB_IN_B16(const_0_16_out),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0F_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0F_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0F_Y09_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0F_Y09_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0F_Y0A_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0F_Y0A_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0F_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0F_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0F_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0F_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0E_Y0A_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0E_Y0A_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0F_Y0A_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0F_Y0A_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(const_0_1_out),
    .SB_T1_EAST_SB_IN_B16(const_0_16_out),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0F_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0F_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0F_Y09_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0F_Y09_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0F_Y0A_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0F_Y0A_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0F_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0F_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0F_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0F_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0E_Y0A_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0E_Y0A_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0F_Y0A_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0F_Y0A_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(const_0_1_out),
    .SB_T2_EAST_SB_IN_B16(const_0_16_out),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0F_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0F_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0F_Y09_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0F_Y09_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0F_Y0A_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0F_Y0A_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0F_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0F_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0F_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0F_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0E_Y0A_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0E_Y0A_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0F_Y0A_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0F_Y0A_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(const_0_1_out),
    .SB_T3_EAST_SB_IN_B16(const_0_16_out),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0F_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0F_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0F_Y09_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0F_Y09_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0F_Y0A_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0F_Y0A_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0F_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0F_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0F_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0F_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0E_Y0A_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0E_Y0A_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0F_Y0A_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0F_Y0A_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(const_0_1_out),
    .SB_T4_EAST_SB_IN_B16(const_0_16_out),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0F_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0F_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0F_Y09_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0F_Y09_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0F_Y0A_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0F_Y0A_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0F_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0F_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0F_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0F_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0E_Y0A_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0E_Y0A_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0F_Y0A_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0F_Y0A_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y0A_clk_pass_through_out_right),
    .clk_out(Tile_X0F_Y0A_clk_out),
    .config_config_addr(Tile_X0F_Y09_config_out_config_addr),
    .config_config_data(Tile_X0F_Y09_config_out_config_data),
    .config_out_config_addr(Tile_X0F_Y0A_config_out_config_addr),
    .config_out_config_data(Tile_X0F_Y0A_config_out_config_data),
    .config_out_read(Tile_X0F_Y0A_config_out_read),
    .config_out_write(Tile_X0F_Y0A_config_out_write),
    .config_read(Tile_X0F_Y09_config_out_read),
    .config_write(Tile_X0F_Y09_config_out_write),
    .hi(Tile_X0F_Y0A_hi_unq1),
    .lo(Tile_X0F_Y0A_lo_unq1),
    .read_config_data(Tile_X0F_Y0A_read_config_data),
    .read_config_data_in(Tile_X0F_Y09_read_config_data),
    .reset(Tile_X0F_Y09_reset_out),
    .reset_out(Tile_X0F_Y0A_reset_out),
    .stall(Tile_X0F_Y09_stall_out),
    .stall_out(Tile_X0F_Y0A_stall_out),
    .tile_id(Tile_X0F_Y0A_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0F_Y0A_hi (
    .in(Tile_X0F_Y0A_hi_unq1),
    .out(Tile_X0F_Y0A_hi_out)
);
mantle_wire__typeBit8 Tile_X0F_Y0A_lo (
    .in(Tile_X0F_Y0A_lo_unq1),
    .out(Tile_X0F_Y0A_lo_out)
);
wire [15:0] Tile_X0F_Y0A_tile_id_out;
assign Tile_X0F_Y0A_tile_id_out = {Tile_X0F_Y0A_lo_out[7],Tile_X0F_Y0A_lo_out[7:6],Tile_X0F_Y0A_lo_out[6],Tile_X0F_Y0A_hi_out[6:5],Tile_X0F_Y0A_hi_out[5:4],Tile_X0F_Y0A_lo_out[3],Tile_X0F_Y0A_lo_out[3:2],Tile_X0F_Y0A_lo_out[2],Tile_X0F_Y0A_hi_out[2],Tile_X0F_Y0A_lo_out[1],Tile_X0F_Y0A_hi_out[1],Tile_X0F_Y0A_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0F_Y0A_tile_id (
    .in(Tile_X0F_Y0A_tile_id_in),
    .out(Tile_X0F_Y0A_tile_id_out)
);
Tile_MemCore Tile_X0F_Y0B (
    .SB_T0_EAST_SB_IN_B1(const_0_1_out),
    .SB_T0_EAST_SB_IN_B16(const_0_16_out),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0F_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0F_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0F_Y0A_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0F_Y0A_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0F_Y0B_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0F_Y0B_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0F_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0F_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0F_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0F_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0E_Y0B_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0E_Y0B_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0F_Y0B_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0F_Y0B_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(const_0_1_out),
    .SB_T1_EAST_SB_IN_B16(const_0_16_out),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0F_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0F_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0F_Y0A_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0F_Y0A_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0F_Y0B_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0F_Y0B_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0F_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0F_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0F_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0F_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0E_Y0B_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0E_Y0B_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0F_Y0B_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0F_Y0B_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(const_0_1_out),
    .SB_T2_EAST_SB_IN_B16(const_0_16_out),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0F_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0F_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0F_Y0A_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0F_Y0A_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0F_Y0B_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0F_Y0B_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0F_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0F_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0F_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0F_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0E_Y0B_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0E_Y0B_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0F_Y0B_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0F_Y0B_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(const_0_1_out),
    .SB_T3_EAST_SB_IN_B16(const_0_16_out),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0F_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0F_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0F_Y0A_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0F_Y0A_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0F_Y0B_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0F_Y0B_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0F_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0F_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0F_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0F_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0E_Y0B_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0E_Y0B_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0F_Y0B_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0F_Y0B_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(const_0_1_out),
    .SB_T4_EAST_SB_IN_B16(const_0_16_out),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0F_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0F_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0F_Y0A_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0F_Y0A_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0F_Y0B_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0F_Y0B_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0F_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0F_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0F_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0F_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0E_Y0B_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0E_Y0B_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0F_Y0B_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0F_Y0B_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y0B_clk_pass_through_out_right),
    .clk_out(Tile_X0F_Y0B_clk_out),
    .config_config_addr(Tile_X0F_Y0A_config_out_config_addr),
    .config_config_data(Tile_X0F_Y0A_config_out_config_data),
    .config_out_config_addr(Tile_X0F_Y0B_config_out_config_addr),
    .config_out_config_data(Tile_X0F_Y0B_config_out_config_data),
    .config_out_read(Tile_X0F_Y0B_config_out_read),
    .config_out_write(Tile_X0F_Y0B_config_out_write),
    .config_read(Tile_X0F_Y0A_config_out_read),
    .config_write(Tile_X0F_Y0A_config_out_write),
    .hi(Tile_X0F_Y0B_hi_unq1),
    .lo(Tile_X0F_Y0B_lo_unq1),
    .read_config_data(Tile_X0F_Y0B_read_config_data),
    .read_config_data_in(Tile_X0F_Y0A_read_config_data),
    .reset(Tile_X0F_Y0A_reset_out),
    .reset_out(Tile_X0F_Y0B_reset_out),
    .stall(Tile_X0F_Y0A_stall_out),
    .stall_out(Tile_X0F_Y0B_stall_out),
    .tile_id(Tile_X0F_Y0B_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0F_Y0B_hi (
    .in(Tile_X0F_Y0B_hi_unq1),
    .out(Tile_X0F_Y0B_hi_out)
);
mantle_wire__typeBit8 Tile_X0F_Y0B_lo (
    .in(Tile_X0F_Y0B_lo_unq1),
    .out(Tile_X0F_Y0B_lo_out)
);
wire [15:0] Tile_X0F_Y0B_tile_id_out;
assign Tile_X0F_Y0B_tile_id_out = {Tile_X0F_Y0B_lo_out[7],Tile_X0F_Y0B_lo_out[7:6],Tile_X0F_Y0B_lo_out[6],Tile_X0F_Y0B_hi_out[6:5],Tile_X0F_Y0B_hi_out[5:4],Tile_X0F_Y0B_lo_out[3],Tile_X0F_Y0B_lo_out[3:2],Tile_X0F_Y0B_lo_out[2],Tile_X0F_Y0B_hi_out[2],Tile_X0F_Y0B_lo_out[1],Tile_X0F_Y0B_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X0F_Y0B_tile_id (
    .in(Tile_X0F_Y0B_tile_id_in),
    .out(Tile_X0F_Y0B_tile_id_out)
);
Tile_MemCore Tile_X0F_Y0C (
    .SB_T0_EAST_SB_IN_B1(const_0_1_out),
    .SB_T0_EAST_SB_IN_B16(const_0_16_out),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0F_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0F_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0F_Y0B_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0F_Y0B_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0F_Y0C_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0F_Y0C_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0F_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0F_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0F_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0F_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0E_Y0C_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0E_Y0C_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0F_Y0C_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0F_Y0C_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(const_0_1_out),
    .SB_T1_EAST_SB_IN_B16(const_0_16_out),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0F_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0F_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0F_Y0B_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0F_Y0B_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0F_Y0C_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0F_Y0C_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0F_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0F_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0F_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0F_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0E_Y0C_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0E_Y0C_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0F_Y0C_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0F_Y0C_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(const_0_1_out),
    .SB_T2_EAST_SB_IN_B16(const_0_16_out),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0F_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0F_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0F_Y0B_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0F_Y0B_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0F_Y0C_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0F_Y0C_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0F_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0F_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0F_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0F_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0E_Y0C_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0E_Y0C_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0F_Y0C_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0F_Y0C_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(const_0_1_out),
    .SB_T3_EAST_SB_IN_B16(const_0_16_out),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0F_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0F_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0F_Y0B_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0F_Y0B_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0F_Y0C_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0F_Y0C_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0F_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0F_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0F_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0F_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0E_Y0C_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0E_Y0C_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0F_Y0C_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0F_Y0C_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(const_0_1_out),
    .SB_T4_EAST_SB_IN_B16(const_0_16_out),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0F_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0F_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0F_Y0B_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0F_Y0B_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0F_Y0C_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0F_Y0C_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0F_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0F_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0F_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0F_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0E_Y0C_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0E_Y0C_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0F_Y0C_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0F_Y0C_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y0C_clk_pass_through_out_right),
    .clk_out(Tile_X0F_Y0C_clk_out),
    .config_config_addr(Tile_X0F_Y0B_config_out_config_addr),
    .config_config_data(Tile_X0F_Y0B_config_out_config_data),
    .config_out_config_addr(Tile_X0F_Y0C_config_out_config_addr),
    .config_out_config_data(Tile_X0F_Y0C_config_out_config_data),
    .config_out_read(Tile_X0F_Y0C_config_out_read),
    .config_out_write(Tile_X0F_Y0C_config_out_write),
    .config_read(Tile_X0F_Y0B_config_out_read),
    .config_write(Tile_X0F_Y0B_config_out_write),
    .hi(Tile_X0F_Y0C_hi_unq1),
    .lo(Tile_X0F_Y0C_lo_unq1),
    .read_config_data(Tile_X0F_Y0C_read_config_data),
    .read_config_data_in(Tile_X0F_Y0B_read_config_data),
    .reset(Tile_X0F_Y0B_reset_out),
    .reset_out(Tile_X0F_Y0C_reset_out),
    .stall(Tile_X0F_Y0B_stall_out),
    .stall_out(Tile_X0F_Y0C_stall_out),
    .tile_id(Tile_X0F_Y0C_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0F_Y0C_hi (
    .in(Tile_X0F_Y0C_hi_unq1),
    .out(Tile_X0F_Y0C_hi_out)
);
mantle_wire__typeBit8 Tile_X0F_Y0C_lo (
    .in(Tile_X0F_Y0C_lo_unq1),
    .out(Tile_X0F_Y0C_lo_out)
);
wire [15:0] Tile_X0F_Y0C_tile_id_out;
assign Tile_X0F_Y0C_tile_id_out = {Tile_X0F_Y0C_lo_out[7],Tile_X0F_Y0C_lo_out[7:6],Tile_X0F_Y0C_lo_out[6],Tile_X0F_Y0C_hi_out[6:5],Tile_X0F_Y0C_hi_out[5:4],Tile_X0F_Y0C_lo_out[3],Tile_X0F_Y0C_lo_out[3:2],Tile_X0F_Y0C_lo_out[2],Tile_X0F_Y0C_hi_out[2:1],Tile_X0F_Y0C_lo_out[0],Tile_X0F_Y0C_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0F_Y0C_tile_id (
    .in(Tile_X0F_Y0C_tile_id_in),
    .out(Tile_X0F_Y0C_tile_id_out)
);
Tile_MemCore Tile_X0F_Y0D (
    .SB_T0_EAST_SB_IN_B1(const_0_1_out),
    .SB_T0_EAST_SB_IN_B16(const_0_16_out),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0F_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0F_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0F_Y0C_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0F_Y0C_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0F_Y0D_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0F_Y0D_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0F_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0F_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0F_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0F_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0E_Y0D_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0E_Y0D_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0F_Y0D_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0F_Y0D_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(const_0_1_out),
    .SB_T1_EAST_SB_IN_B16(const_0_16_out),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0F_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0F_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0F_Y0C_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0F_Y0C_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0F_Y0D_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0F_Y0D_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0F_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0F_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0F_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0F_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0E_Y0D_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0E_Y0D_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0F_Y0D_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0F_Y0D_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(const_0_1_out),
    .SB_T2_EAST_SB_IN_B16(const_0_16_out),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0F_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0F_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0F_Y0C_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0F_Y0C_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0F_Y0D_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0F_Y0D_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0F_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0F_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0F_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0F_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0E_Y0D_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0E_Y0D_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0F_Y0D_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0F_Y0D_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(const_0_1_out),
    .SB_T3_EAST_SB_IN_B16(const_0_16_out),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0F_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0F_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0F_Y0C_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0F_Y0C_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0F_Y0D_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0F_Y0D_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0F_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0F_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0F_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0F_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0E_Y0D_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0E_Y0D_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0F_Y0D_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0F_Y0D_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(const_0_1_out),
    .SB_T4_EAST_SB_IN_B16(const_0_16_out),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0F_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0F_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0F_Y0C_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0F_Y0C_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0F_Y0D_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0F_Y0D_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0F_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0F_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0F_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0F_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0E_Y0D_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0E_Y0D_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0F_Y0D_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0F_Y0D_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y0D_clk_pass_through_out_right),
    .clk_out(Tile_X0F_Y0D_clk_out),
    .config_config_addr(Tile_X0F_Y0C_config_out_config_addr),
    .config_config_data(Tile_X0F_Y0C_config_out_config_data),
    .config_out_config_addr(Tile_X0F_Y0D_config_out_config_addr),
    .config_out_config_data(Tile_X0F_Y0D_config_out_config_data),
    .config_out_read(Tile_X0F_Y0D_config_out_read),
    .config_out_write(Tile_X0F_Y0D_config_out_write),
    .config_read(Tile_X0F_Y0C_config_out_read),
    .config_write(Tile_X0F_Y0C_config_out_write),
    .hi(Tile_X0F_Y0D_hi_unq1),
    .lo(Tile_X0F_Y0D_lo_unq1),
    .read_config_data(Tile_X0F_Y0D_read_config_data),
    .read_config_data_in(Tile_X0F_Y0C_read_config_data),
    .reset(Tile_X0F_Y0C_reset_out),
    .reset_out(Tile_X0F_Y0D_reset_out),
    .stall(Tile_X0F_Y0C_stall_out),
    .stall_out(Tile_X0F_Y0D_stall_out),
    .tile_id(Tile_X0F_Y0D_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0F_Y0D_hi (
    .in(Tile_X0F_Y0D_hi_unq1),
    .out(Tile_X0F_Y0D_hi_out)
);
mantle_wire__typeBit8 Tile_X0F_Y0D_lo (
    .in(Tile_X0F_Y0D_lo_unq1),
    .out(Tile_X0F_Y0D_lo_out)
);
wire [15:0] Tile_X0F_Y0D_tile_id_out;
assign Tile_X0F_Y0D_tile_id_out = {Tile_X0F_Y0D_lo_out[7],Tile_X0F_Y0D_lo_out[7:6],Tile_X0F_Y0D_lo_out[6],Tile_X0F_Y0D_hi_out[6:5],Tile_X0F_Y0D_hi_out[5:4],Tile_X0F_Y0D_lo_out[3],Tile_X0F_Y0D_lo_out[3:2],Tile_X0F_Y0D_lo_out[2],Tile_X0F_Y0D_hi_out[2:1],Tile_X0F_Y0D_lo_out[0],Tile_X0F_Y0D_hi_out[0]};
mantle_wire__typeBitIn16 Tile_X0F_Y0D_tile_id (
    .in(Tile_X0F_Y0D_tile_id_in),
    .out(Tile_X0F_Y0D_tile_id_out)
);
Tile_MemCore Tile_X0F_Y0E (
    .SB_T0_EAST_SB_IN_B1(const_0_1_out),
    .SB_T0_EAST_SB_IN_B16(const_0_16_out),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0F_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0F_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0F_Y0D_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0F_Y0D_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0F_Y0E_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0F_Y0E_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0F_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0F_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0F_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0F_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0E_Y0E_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0E_Y0E_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0F_Y0E_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0F_Y0E_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(const_0_1_out),
    .SB_T1_EAST_SB_IN_B16(const_0_16_out),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0F_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0F_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0F_Y0D_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0F_Y0D_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0F_Y0E_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0F_Y0E_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0F_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0F_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0F_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0F_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0E_Y0E_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0E_Y0E_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0F_Y0E_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0F_Y0E_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(const_0_1_out),
    .SB_T2_EAST_SB_IN_B16(const_0_16_out),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0F_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0F_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0F_Y0D_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0F_Y0D_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0F_Y0E_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0F_Y0E_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0F_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0F_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0F_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0F_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0E_Y0E_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0E_Y0E_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0F_Y0E_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0F_Y0E_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(const_0_1_out),
    .SB_T3_EAST_SB_IN_B16(const_0_16_out),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0F_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0F_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0F_Y0D_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0F_Y0D_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0F_Y0E_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0F_Y0E_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0F_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0F_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0F_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0F_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0E_Y0E_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0E_Y0E_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0F_Y0E_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0F_Y0E_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(const_0_1_out),
    .SB_T4_EAST_SB_IN_B16(const_0_16_out),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0F_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0F_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0F_Y0D_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0F_Y0D_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0F_Y0E_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0F_Y0E_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0F_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0F_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0F_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0F_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0E_Y0E_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0E_Y0E_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0F_Y0E_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0F_Y0E_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y0E_clk_pass_through_out_right),
    .clk_out(Tile_X0F_Y0E_clk_out),
    .config_config_addr(Tile_X0F_Y0D_config_out_config_addr),
    .config_config_data(Tile_X0F_Y0D_config_out_config_data),
    .config_out_config_addr(Tile_X0F_Y0E_config_out_config_addr),
    .config_out_config_data(Tile_X0F_Y0E_config_out_config_data),
    .config_out_read(Tile_X0F_Y0E_config_out_read),
    .config_out_write(Tile_X0F_Y0E_config_out_write),
    .config_read(Tile_X0F_Y0D_config_out_read),
    .config_write(Tile_X0F_Y0D_config_out_write),
    .hi(Tile_X0F_Y0E_hi_unq1),
    .lo(Tile_X0F_Y0E_lo_unq1),
    .read_config_data(Tile_X0F_Y0E_read_config_data),
    .read_config_data_in(Tile_X0F_Y0D_read_config_data),
    .reset(Tile_X0F_Y0D_reset_out),
    .reset_out(Tile_X0F_Y0E_reset_out),
    .stall(Tile_X0F_Y0D_stall_out),
    .stall_out(Tile_X0F_Y0E_stall_out),
    .tile_id(Tile_X0F_Y0E_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0F_Y0E_hi (
    .in(Tile_X0F_Y0E_hi_unq1),
    .out(Tile_X0F_Y0E_hi_out)
);
mantle_wire__typeBit8 Tile_X0F_Y0E_lo (
    .in(Tile_X0F_Y0E_lo_unq1),
    .out(Tile_X0F_Y0E_lo_out)
);
wire [15:0] Tile_X0F_Y0E_tile_id_out;
assign Tile_X0F_Y0E_tile_id_out = {Tile_X0F_Y0E_lo_out[7],Tile_X0F_Y0E_lo_out[7:6],Tile_X0F_Y0E_lo_out[6],Tile_X0F_Y0E_hi_out[6:5],Tile_X0F_Y0E_hi_out[5:4],Tile_X0F_Y0E_lo_out[3],Tile_X0F_Y0E_lo_out[3:2],Tile_X0F_Y0E_lo_out[2],Tile_X0F_Y0E_hi_out[2:1],Tile_X0F_Y0E_hi_out[1],Tile_X0F_Y0E_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0F_Y0E_tile_id (
    .in(Tile_X0F_Y0E_tile_id_in),
    .out(Tile_X0F_Y0E_tile_id_out)
);
Tile_MemCore Tile_X0F_Y0F (
    .SB_T0_EAST_SB_IN_B1(const_0_1_out),
    .SB_T0_EAST_SB_IN_B16(const_0_16_out),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0F_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0F_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0F_Y0E_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0F_Y0E_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0F_Y0F_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0F_Y0F_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(Tile_X0F_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_IN_B16(Tile_X0F_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0F_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0F_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0E_Y0F_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0E_Y0F_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0F_Y0F_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0F_Y0F_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(const_0_1_out),
    .SB_T1_EAST_SB_IN_B16(const_0_16_out),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0F_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0F_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0F_Y0E_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0F_Y0E_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0F_Y0F_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0F_Y0F_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(Tile_X0F_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_IN_B16(Tile_X0F_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0F_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0F_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0E_Y0F_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0E_Y0F_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0F_Y0F_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0F_Y0F_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(const_0_1_out),
    .SB_T2_EAST_SB_IN_B16(const_0_16_out),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0F_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0F_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0F_Y0E_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0F_Y0E_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0F_Y0F_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0F_Y0F_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(Tile_X0F_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_IN_B16(Tile_X0F_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0F_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0F_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0E_Y0F_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0E_Y0F_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0F_Y0F_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0F_Y0F_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(const_0_1_out),
    .SB_T3_EAST_SB_IN_B16(const_0_16_out),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0F_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0F_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0F_Y0E_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0F_Y0E_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0F_Y0F_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0F_Y0F_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(Tile_X0F_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_IN_B16(Tile_X0F_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0F_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0F_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0E_Y0F_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0E_Y0F_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0F_Y0F_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0F_Y0F_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(const_0_1_out),
    .SB_T4_EAST_SB_IN_B16(const_0_16_out),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0F_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0F_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0F_Y0E_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0F_Y0E_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0F_Y0F_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0F_Y0F_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(Tile_X0F_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_IN_B16(Tile_X0F_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0F_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0F_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0E_Y0F_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0E_Y0F_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0F_Y0F_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0F_Y0F_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y0F_clk_pass_through_out_right),
    .clk_out(Tile_X0F_Y0F_clk_out),
    .config_config_addr(Tile_X0F_Y0E_config_out_config_addr),
    .config_config_data(Tile_X0F_Y0E_config_out_config_data),
    .config_out_config_addr(Tile_X0F_Y0F_config_out_config_addr),
    .config_out_config_data(Tile_X0F_Y0F_config_out_config_data),
    .config_out_read(Tile_X0F_Y0F_config_out_read),
    .config_out_write(Tile_X0F_Y0F_config_out_write),
    .config_read(Tile_X0F_Y0E_config_out_read),
    .config_write(Tile_X0F_Y0E_config_out_write),
    .hi(Tile_X0F_Y0F_hi_unq1),
    .lo(Tile_X0F_Y0F_lo_unq1),
    .read_config_data(Tile_X0F_Y0F_read_config_data),
    .read_config_data_in(Tile_X0F_Y0E_read_config_data),
    .reset(Tile_X0F_Y0E_reset_out),
    .reset_out(Tile_X0F_Y0F_reset_out),
    .stall(Tile_X0F_Y0E_stall_out),
    .stall_out(Tile_X0F_Y0F_stall_out),
    .tile_id(Tile_X0F_Y0F_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0F_Y0F_hi (
    .in(Tile_X0F_Y0F_hi_unq1),
    .out(Tile_X0F_Y0F_hi_out)
);
mantle_wire__typeBit8 Tile_X0F_Y0F_lo (
    .in(Tile_X0F_Y0F_lo_unq1),
    .out(Tile_X0F_Y0F_lo_out)
);
wire [15:0] Tile_X0F_Y0F_tile_id_out;
assign Tile_X0F_Y0F_tile_id_out = {Tile_X0F_Y0F_lo_out[7],Tile_X0F_Y0F_lo_out[7:6],Tile_X0F_Y0F_lo_out[6],Tile_X0F_Y0F_hi_out[6:5],Tile_X0F_Y0F_hi_out[5:4],Tile_X0F_Y0F_lo_out[3],Tile_X0F_Y0F_lo_out[3:2],Tile_X0F_Y0F_lo_out[2],Tile_X0F_Y0F_hi_out[2:1],Tile_X0F_Y0F_hi_out[1:0]};
mantle_wire__typeBitIn16 Tile_X0F_Y0F_tile_id (
    .in(Tile_X0F_Y0F_tile_id_in),
    .out(Tile_X0F_Y0F_tile_id_out)
);
Tile_MemCore Tile_X0F_Y10 (
    .SB_T0_EAST_SB_IN_B1(const_0_1_out),
    .SB_T0_EAST_SB_IN_B16(const_0_16_out),
    .SB_T0_EAST_SB_OUT_B1(Tile_X0F_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_EAST_SB_OUT_B16(Tile_X0F_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_NORTH_SB_IN_B1(Tile_X0F_Y0F_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_IN_B16(Tile_X0F_Y0F_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_NORTH_SB_OUT_B1(Tile_X0F_Y10_SB_T0_NORTH_SB_OUT_B1),
    .SB_T0_NORTH_SB_OUT_B16(Tile_X0F_Y10_SB_T0_NORTH_SB_OUT_B16),
    .SB_T0_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T0_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T0_SOUTH_SB_OUT_B1(Tile_X0F_Y10_SB_T0_SOUTH_SB_OUT_B1),
    .SB_T0_SOUTH_SB_OUT_B16(Tile_X0F_Y10_SB_T0_SOUTH_SB_OUT_B16),
    .SB_T0_WEST_SB_IN_B1(Tile_X0E_Y10_SB_T0_EAST_SB_OUT_B1),
    .SB_T0_WEST_SB_IN_B16(Tile_X0E_Y10_SB_T0_EAST_SB_OUT_B16),
    .SB_T0_WEST_SB_OUT_B1(Tile_X0F_Y10_SB_T0_WEST_SB_OUT_B1),
    .SB_T0_WEST_SB_OUT_B16(Tile_X0F_Y10_SB_T0_WEST_SB_OUT_B16),
    .SB_T1_EAST_SB_IN_B1(const_0_1_out),
    .SB_T1_EAST_SB_IN_B16(const_0_16_out),
    .SB_T1_EAST_SB_OUT_B1(Tile_X0F_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_EAST_SB_OUT_B16(Tile_X0F_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_NORTH_SB_IN_B1(Tile_X0F_Y0F_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_IN_B16(Tile_X0F_Y0F_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_NORTH_SB_OUT_B1(Tile_X0F_Y10_SB_T1_NORTH_SB_OUT_B1),
    .SB_T1_NORTH_SB_OUT_B16(Tile_X0F_Y10_SB_T1_NORTH_SB_OUT_B16),
    .SB_T1_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T1_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T1_SOUTH_SB_OUT_B1(Tile_X0F_Y10_SB_T1_SOUTH_SB_OUT_B1),
    .SB_T1_SOUTH_SB_OUT_B16(Tile_X0F_Y10_SB_T1_SOUTH_SB_OUT_B16),
    .SB_T1_WEST_SB_IN_B1(Tile_X0E_Y10_SB_T1_EAST_SB_OUT_B1),
    .SB_T1_WEST_SB_IN_B16(Tile_X0E_Y10_SB_T1_EAST_SB_OUT_B16),
    .SB_T1_WEST_SB_OUT_B1(Tile_X0F_Y10_SB_T1_WEST_SB_OUT_B1),
    .SB_T1_WEST_SB_OUT_B16(Tile_X0F_Y10_SB_T1_WEST_SB_OUT_B16),
    .SB_T2_EAST_SB_IN_B1(const_0_1_out),
    .SB_T2_EAST_SB_IN_B16(const_0_16_out),
    .SB_T2_EAST_SB_OUT_B1(Tile_X0F_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_EAST_SB_OUT_B16(Tile_X0F_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_NORTH_SB_IN_B1(Tile_X0F_Y0F_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_IN_B16(Tile_X0F_Y0F_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_NORTH_SB_OUT_B1(Tile_X0F_Y10_SB_T2_NORTH_SB_OUT_B1),
    .SB_T2_NORTH_SB_OUT_B16(Tile_X0F_Y10_SB_T2_NORTH_SB_OUT_B16),
    .SB_T2_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T2_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T2_SOUTH_SB_OUT_B1(Tile_X0F_Y10_SB_T2_SOUTH_SB_OUT_B1),
    .SB_T2_SOUTH_SB_OUT_B16(Tile_X0F_Y10_SB_T2_SOUTH_SB_OUT_B16),
    .SB_T2_WEST_SB_IN_B1(Tile_X0E_Y10_SB_T2_EAST_SB_OUT_B1),
    .SB_T2_WEST_SB_IN_B16(Tile_X0E_Y10_SB_T2_EAST_SB_OUT_B16),
    .SB_T2_WEST_SB_OUT_B1(Tile_X0F_Y10_SB_T2_WEST_SB_OUT_B1),
    .SB_T2_WEST_SB_OUT_B16(Tile_X0F_Y10_SB_T2_WEST_SB_OUT_B16),
    .SB_T3_EAST_SB_IN_B1(const_0_1_out),
    .SB_T3_EAST_SB_IN_B16(const_0_16_out),
    .SB_T3_EAST_SB_OUT_B1(Tile_X0F_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_EAST_SB_OUT_B16(Tile_X0F_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_NORTH_SB_IN_B1(Tile_X0F_Y0F_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_IN_B16(Tile_X0F_Y0F_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_NORTH_SB_OUT_B1(Tile_X0F_Y10_SB_T3_NORTH_SB_OUT_B1),
    .SB_T3_NORTH_SB_OUT_B16(Tile_X0F_Y10_SB_T3_NORTH_SB_OUT_B16),
    .SB_T3_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T3_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T3_SOUTH_SB_OUT_B1(Tile_X0F_Y10_SB_T3_SOUTH_SB_OUT_B1),
    .SB_T3_SOUTH_SB_OUT_B16(Tile_X0F_Y10_SB_T3_SOUTH_SB_OUT_B16),
    .SB_T3_WEST_SB_IN_B1(Tile_X0E_Y10_SB_T3_EAST_SB_OUT_B1),
    .SB_T3_WEST_SB_IN_B16(Tile_X0E_Y10_SB_T3_EAST_SB_OUT_B16),
    .SB_T3_WEST_SB_OUT_B1(Tile_X0F_Y10_SB_T3_WEST_SB_OUT_B1),
    .SB_T3_WEST_SB_OUT_B16(Tile_X0F_Y10_SB_T3_WEST_SB_OUT_B16),
    .SB_T4_EAST_SB_IN_B1(const_0_1_out),
    .SB_T4_EAST_SB_IN_B16(const_0_16_out),
    .SB_T4_EAST_SB_OUT_B1(Tile_X0F_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_EAST_SB_OUT_B16(Tile_X0F_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_NORTH_SB_IN_B1(Tile_X0F_Y0F_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_IN_B16(Tile_X0F_Y0F_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_NORTH_SB_OUT_B1(Tile_X0F_Y10_SB_T4_NORTH_SB_OUT_B1),
    .SB_T4_NORTH_SB_OUT_B16(Tile_X0F_Y10_SB_T4_NORTH_SB_OUT_B16),
    .SB_T4_SOUTH_SB_IN_B1(const_0_1_out),
    .SB_T4_SOUTH_SB_IN_B16(const_0_16_out),
    .SB_T4_SOUTH_SB_OUT_B1(Tile_X0F_Y10_SB_T4_SOUTH_SB_OUT_B1),
    .SB_T4_SOUTH_SB_OUT_B16(Tile_X0F_Y10_SB_T4_SOUTH_SB_OUT_B16),
    .SB_T4_WEST_SB_IN_B1(Tile_X0E_Y10_SB_T4_EAST_SB_OUT_B1),
    .SB_T4_WEST_SB_IN_B16(Tile_X0E_Y10_SB_T4_EAST_SB_OUT_B16),
    .SB_T4_WEST_SB_OUT_B1(Tile_X0F_Y10_SB_T4_WEST_SB_OUT_B1),
    .SB_T4_WEST_SB_OUT_B16(Tile_X0F_Y10_SB_T4_WEST_SB_OUT_B16),
    .clk(Tile_X0E_Y10_clk_pass_through_out_right),
    .clk_out(Tile_X0F_Y10_clk_out),
    .config_config_addr(Tile_X0F_Y0F_config_out_config_addr),
    .config_config_data(Tile_X0F_Y0F_config_out_config_data),
    .config_out_config_addr(Tile_X0F_Y10_config_out_config_addr),
    .config_out_config_data(Tile_X0F_Y10_config_out_config_data),
    .config_out_read(Tile_X0F_Y10_config_out_read),
    .config_out_write(Tile_X0F_Y10_config_out_write),
    .config_read(Tile_X0F_Y0F_config_out_read),
    .config_write(Tile_X0F_Y0F_config_out_write),
    .hi(Tile_X0F_Y10_hi_unq1),
    .lo(Tile_X0F_Y10_lo_unq1),
    .read_config_data(Tile_X0F_Y10_read_config_data),
    .read_config_data_in(Tile_X0F_Y0F_read_config_data),
    .reset(Tile_X0F_Y0F_reset_out),
    .reset_out(Tile_X0F_Y10_reset_out),
    .stall(Tile_X0F_Y0F_stall_out),
    .stall_out(Tile_X0F_Y10_stall_out),
    .tile_id(Tile_X0F_Y10_tile_id_in)
);
mantle_wire__typeBit9 Tile_X0F_Y10_hi (
    .in(Tile_X0F_Y10_hi_unq1),
    .out(Tile_X0F_Y10_hi_out)
);
mantle_wire__typeBit8 Tile_X0F_Y10_lo (
    .in(Tile_X0F_Y10_lo_unq1),
    .out(Tile_X0F_Y10_lo_out)
);
wire [15:0] Tile_X0F_Y10_tile_id_out;
assign Tile_X0F_Y10_tile_id_out = {Tile_X0F_Y10_lo_out[7],Tile_X0F_Y10_lo_out[7:6],Tile_X0F_Y10_lo_out[6],Tile_X0F_Y10_hi_out[6:5],Tile_X0F_Y10_hi_out[5:4],Tile_X0F_Y10_lo_out[3],Tile_X0F_Y10_lo_out[3:2],Tile_X0F_Y10_hi_out[2],Tile_X0F_Y10_lo_out[1],Tile_X0F_Y10_lo_out[1:0],Tile_X0F_Y10_lo_out[0]};
mantle_wire__typeBitIn16 Tile_X0F_Y10_tile_id (
    .in(Tile_X0F_Y10_tile_id_in),
    .out(Tile_X0F_Y10_tile_id_out)
);
coreir_const #(
    .value(1'h0),
    .width(1)
) const_0_1 (
    .out(const_0_1_out)
);
coreir_const #(
    .value(16'h0000),
    .width(16)
) const_0_16 (
    .out(const_0_16_out)
);
coreir_const #(
    .value(32'h00000000),
    .width(32)
) const_0_32 (
    .out(const_0_32_out)
);
Or16x32 read_config_data_or_final (
    .I0(Tile_X00_Y10_read_config_data),
    .I1(Tile_X01_Y10_read_config_data),
    .I2(Tile_X02_Y10_read_config_data),
    .I3(Tile_X03_Y10_read_config_data),
    .I4(Tile_X04_Y10_read_config_data),
    .I5(Tile_X05_Y10_read_config_data),
    .I6(Tile_X06_Y10_read_config_data),
    .I7(Tile_X07_Y10_read_config_data),
    .I8(Tile_X08_Y10_read_config_data),
    .I9(Tile_X09_Y10_read_config_data),
    .I10(Tile_X0A_Y10_read_config_data),
    .I11(Tile_X0B_Y10_read_config_data),
    .I12(Tile_X0C_Y10_read_config_data),
    .I13(Tile_X0D_Y10_read_config_data),
    .I14(Tile_X0E_Y10_read_config_data),
    .I15(Tile_X0F_Y10_read_config_data),
    .O(read_config_data_or_final_O)
);
assign io2glb_16_X00_Y00 = Tile_X00_Y00_io2glb_16;
assign io2glb_16_X01_Y00 = Tile_X01_Y00_io2glb_16;
assign io2glb_16_X02_Y00 = Tile_X02_Y00_io2glb_16;
assign io2glb_16_X03_Y00 = Tile_X03_Y00_io2glb_16;
assign io2glb_16_X04_Y00 = Tile_X04_Y00_io2glb_16;
assign io2glb_16_X05_Y00 = Tile_X05_Y00_io2glb_16;
assign io2glb_16_X06_Y00 = Tile_X06_Y00_io2glb_16;
assign io2glb_16_X07_Y00 = Tile_X07_Y00_io2glb_16;
assign io2glb_16_X08_Y00 = Tile_X08_Y00_io2glb_16;
assign io2glb_16_X09_Y00 = Tile_X09_Y00_io2glb_16;
assign io2glb_16_X0A_Y00 = Tile_X0A_Y00_io2glb_16;
assign io2glb_16_X0B_Y00 = Tile_X0B_Y00_io2glb_16;
assign io2glb_16_X0C_Y00 = Tile_X0C_Y00_io2glb_16;
assign io2glb_16_X0D_Y00 = Tile_X0D_Y00_io2glb_16;
assign io2glb_16_X0E_Y00 = Tile_X0E_Y00_io2glb_16;
assign io2glb_16_X0F_Y00 = Tile_X0F_Y00_io2glb_16;
assign io2glb_1_X00_Y00 = Tile_X00_Y00_io2glb_1;
assign io2glb_1_X01_Y00 = Tile_X01_Y00_io2glb_1;
assign io2glb_1_X02_Y00 = Tile_X02_Y00_io2glb_1;
assign io2glb_1_X03_Y00 = Tile_X03_Y00_io2glb_1;
assign io2glb_1_X04_Y00 = Tile_X04_Y00_io2glb_1;
assign io2glb_1_X05_Y00 = Tile_X05_Y00_io2glb_1;
assign io2glb_1_X06_Y00 = Tile_X06_Y00_io2glb_1;
assign io2glb_1_X07_Y00 = Tile_X07_Y00_io2glb_1;
assign io2glb_1_X08_Y00 = Tile_X08_Y00_io2glb_1;
assign io2glb_1_X09_Y00 = Tile_X09_Y00_io2glb_1;
assign io2glb_1_X0A_Y00 = Tile_X0A_Y00_io2glb_1;
assign io2glb_1_X0B_Y00 = Tile_X0B_Y00_io2glb_1;
assign io2glb_1_X0C_Y00 = Tile_X0C_Y00_io2glb_1;
assign io2glb_1_X0D_Y00 = Tile_X0D_Y00_io2glb_1;
assign io2glb_1_X0E_Y00 = Tile_X0E_Y00_io2glb_1;
assign io2glb_1_X0F_Y00 = Tile_X0F_Y00_io2glb_1;
assign read_config_data = read_config_data_or_final_O;
endmodule

module Garnet (
    input clk,
    input [31:0] config_0_config_addr,
    input [31:0] config_0_config_data,
    input [0:0] config_0_read,
    input [0:0] config_0_write,
    input [31:0] config_10_config_addr,
    input [31:0] config_10_config_data,
    input [0:0] config_10_read,
    input [0:0] config_10_write,
    input [31:0] config_11_config_addr,
    input [31:0] config_11_config_data,
    input [0:0] config_11_read,
    input [0:0] config_11_write,
    input [31:0] config_12_config_addr,
    input [31:0] config_12_config_data,
    input [0:0] config_12_read,
    input [0:0] config_12_write,
    input [31:0] config_13_config_addr,
    input [31:0] config_13_config_data,
    input [0:0] config_13_read,
    input [0:0] config_13_write,
    input [31:0] config_14_config_addr,
    input [31:0] config_14_config_data,
    input [0:0] config_14_read,
    input [0:0] config_14_write,
    input [31:0] config_15_config_addr,
    input [31:0] config_15_config_data,
    input [0:0] config_15_read,
    input [0:0] config_15_write,
    input [31:0] config_1_config_addr,
    input [31:0] config_1_config_data,
    input [0:0] config_1_read,
    input [0:0] config_1_write,
    input [31:0] config_2_config_addr,
    input [31:0] config_2_config_data,
    input [0:0] config_2_read,
    input [0:0] config_2_write,
    input [31:0] config_3_config_addr,
    input [31:0] config_3_config_data,
    input [0:0] config_3_read,
    input [0:0] config_3_write,
    input [31:0] config_4_config_addr,
    input [31:0] config_4_config_data,
    input [0:0] config_4_read,
    input [0:0] config_4_write,
    input [31:0] config_5_config_addr,
    input [31:0] config_5_config_data,
    input [0:0] config_5_read,
    input [0:0] config_5_write,
    input [31:0] config_6_config_addr,
    input [31:0] config_6_config_data,
    input [0:0] config_6_read,
    input [0:0] config_6_write,
    input [31:0] config_7_config_addr,
    input [31:0] config_7_config_data,
    input [0:0] config_7_read,
    input [0:0] config_7_write,
    input [31:0] config_8_config_addr,
    input [31:0] config_8_config_data,
    input [0:0] config_8_read,
    input [0:0] config_8_write,
    input [31:0] config_9_config_addr,
    input [31:0] config_9_config_data,
    input [0:0] config_9_read,
    input [0:0] config_9_write,
    input [15:0] glb2io_16_X00_Y00,
    input [15:0] glb2io_16_X01_Y00,
    input [15:0] glb2io_16_X02_Y00,
    input [15:0] glb2io_16_X03_Y00,
    input [15:0] glb2io_16_X04_Y00,
    input [15:0] glb2io_16_X05_Y00,
    input [15:0] glb2io_16_X06_Y00,
    input [15:0] glb2io_16_X07_Y00,
    input [15:0] glb2io_16_X08_Y00,
    input [15:0] glb2io_16_X09_Y00,
    input [15:0] glb2io_16_X0A_Y00,
    input [15:0] glb2io_16_X0B_Y00,
    input [15:0] glb2io_16_X0C_Y00,
    input [15:0] glb2io_16_X0D_Y00,
    input [15:0] glb2io_16_X0E_Y00,
    input [15:0] glb2io_16_X0F_Y00,
    input [0:0] glb2io_1_X00_Y00,
    input [0:0] glb2io_1_X01_Y00,
    input [0:0] glb2io_1_X02_Y00,
    input [0:0] glb2io_1_X03_Y00,
    input [0:0] glb2io_1_X04_Y00,
    input [0:0] glb2io_1_X05_Y00,
    input [0:0] glb2io_1_X06_Y00,
    input [0:0] glb2io_1_X07_Y00,
    input [0:0] glb2io_1_X08_Y00,
    input [0:0] glb2io_1_X09_Y00,
    input [0:0] glb2io_1_X0A_Y00,
    input [0:0] glb2io_1_X0B_Y00,
    input [0:0] glb2io_1_X0C_Y00,
    input [0:0] glb2io_1_X0D_Y00,
    input [0:0] glb2io_1_X0E_Y00,
    input [0:0] glb2io_1_X0F_Y00,
    output [15:0] io2glb_16_X00_Y00,
    output [15:0] io2glb_16_X01_Y00,
    output [15:0] io2glb_16_X02_Y00,
    output [15:0] io2glb_16_X03_Y00,
    output [15:0] io2glb_16_X04_Y00,
    output [15:0] io2glb_16_X05_Y00,
    output [15:0] io2glb_16_X06_Y00,
    output [15:0] io2glb_16_X07_Y00,
    output [15:0] io2glb_16_X08_Y00,
    output [15:0] io2glb_16_X09_Y00,
    output [15:0] io2glb_16_X0A_Y00,
    output [15:0] io2glb_16_X0B_Y00,
    output [15:0] io2glb_16_X0C_Y00,
    output [15:0] io2glb_16_X0D_Y00,
    output [15:0] io2glb_16_X0E_Y00,
    output [15:0] io2glb_16_X0F_Y00,
    output [0:0] io2glb_1_X00_Y00,
    output [0:0] io2glb_1_X01_Y00,
    output [0:0] io2glb_1_X02_Y00,
    output [0:0] io2glb_1_X03_Y00,
    output [0:0] io2glb_1_X04_Y00,
    output [0:0] io2glb_1_X05_Y00,
    output [0:0] io2glb_1_X06_Y00,
    output [0:0] io2glb_1_X07_Y00,
    output [0:0] io2glb_1_X08_Y00,
    output [0:0] io2glb_1_X09_Y00,
    output [0:0] io2glb_1_X0A_Y00,
    output [0:0] io2glb_1_X0B_Y00,
    output [0:0] io2glb_1_X0C_Y00,
    output [0:0] io2glb_1_X0D_Y00,
    output [0:0] io2glb_1_X0E_Y00,
    output [0:0] io2glb_1_X0F_Y00,
    output [31:0] read_config_data,
    input reset,
    input [15:0] stall
);
wire [15:0] Interconnect_inst0_io2glb_16_X00_Y00;
wire [15:0] Interconnect_inst0_io2glb_16_X01_Y00;
wire [15:0] Interconnect_inst0_io2glb_16_X02_Y00;
wire [15:0] Interconnect_inst0_io2glb_16_X03_Y00;
wire [15:0] Interconnect_inst0_io2glb_16_X04_Y00;
wire [15:0] Interconnect_inst0_io2glb_16_X05_Y00;
wire [15:0] Interconnect_inst0_io2glb_16_X06_Y00;
wire [15:0] Interconnect_inst0_io2glb_16_X07_Y00;
wire [15:0] Interconnect_inst0_io2glb_16_X08_Y00;
wire [15:0] Interconnect_inst0_io2glb_16_X09_Y00;
wire [15:0] Interconnect_inst0_io2glb_16_X0A_Y00;
wire [15:0] Interconnect_inst0_io2glb_16_X0B_Y00;
wire [15:0] Interconnect_inst0_io2glb_16_X0C_Y00;
wire [15:0] Interconnect_inst0_io2glb_16_X0D_Y00;
wire [15:0] Interconnect_inst0_io2glb_16_X0E_Y00;
wire [15:0] Interconnect_inst0_io2glb_16_X0F_Y00;
wire [0:0] Interconnect_inst0_io2glb_1_X00_Y00;
wire [0:0] Interconnect_inst0_io2glb_1_X01_Y00;
wire [0:0] Interconnect_inst0_io2glb_1_X02_Y00;
wire [0:0] Interconnect_inst0_io2glb_1_X03_Y00;
wire [0:0] Interconnect_inst0_io2glb_1_X04_Y00;
wire [0:0] Interconnect_inst0_io2glb_1_X05_Y00;
wire [0:0] Interconnect_inst0_io2glb_1_X06_Y00;
wire [0:0] Interconnect_inst0_io2glb_1_X07_Y00;
wire [0:0] Interconnect_inst0_io2glb_1_X08_Y00;
wire [0:0] Interconnect_inst0_io2glb_1_X09_Y00;
wire [0:0] Interconnect_inst0_io2glb_1_X0A_Y00;
wire [0:0] Interconnect_inst0_io2glb_1_X0B_Y00;
wire [0:0] Interconnect_inst0_io2glb_1_X0C_Y00;
wire [0:0] Interconnect_inst0_io2glb_1_X0D_Y00;
wire [0:0] Interconnect_inst0_io2glb_1_X0E_Y00;
wire [0:0] Interconnect_inst0_io2glb_1_X0F_Y00;
wire [31:0] Interconnect_inst0_read_config_data;
Interconnect Interconnect_inst0 (
    .clk(clk),
    .config_0_config_addr(config_0_config_addr),
    .config_0_config_data(config_0_config_data),
    .config_0_read(config_0_read),
    .config_0_write(config_0_write),
    .config_10_config_addr(config_10_config_addr),
    .config_10_config_data(config_10_config_data),
    .config_10_read(config_10_read),
    .config_10_write(config_10_write),
    .config_11_config_addr(config_11_config_addr),
    .config_11_config_data(config_11_config_data),
    .config_11_read(config_11_read),
    .config_11_write(config_11_write),
    .config_12_config_addr(config_12_config_addr),
    .config_12_config_data(config_12_config_data),
    .config_12_read(config_12_read),
    .config_12_write(config_12_write),
    .config_13_config_addr(config_13_config_addr),
    .config_13_config_data(config_13_config_data),
    .config_13_read(config_13_read),
    .config_13_write(config_13_write),
    .config_14_config_addr(config_14_config_addr),
    .config_14_config_data(config_14_config_data),
    .config_14_read(config_14_read),
    .config_14_write(config_14_write),
    .config_15_config_addr(config_15_config_addr),
    .config_15_config_data(config_15_config_data),
    .config_15_read(config_15_read),
    .config_15_write(config_15_write),
    .config_1_config_addr(config_1_config_addr),
    .config_1_config_data(config_1_config_data),
    .config_1_read(config_1_read),
    .config_1_write(config_1_write),
    .config_2_config_addr(config_2_config_addr),
    .config_2_config_data(config_2_config_data),
    .config_2_read(config_2_read),
    .config_2_write(config_2_write),
    .config_3_config_addr(config_3_config_addr),
    .config_3_config_data(config_3_config_data),
    .config_3_read(config_3_read),
    .config_3_write(config_3_write),
    .config_4_config_addr(config_4_config_addr),
    .config_4_config_data(config_4_config_data),
    .config_4_read(config_4_read),
    .config_4_write(config_4_write),
    .config_5_config_addr(config_5_config_addr),
    .config_5_config_data(config_5_config_data),
    .config_5_read(config_5_read),
    .config_5_write(config_5_write),
    .config_6_config_addr(config_6_config_addr),
    .config_6_config_data(config_6_config_data),
    .config_6_read(config_6_read),
    .config_6_write(config_6_write),
    .config_7_config_addr(config_7_config_addr),
    .config_7_config_data(config_7_config_data),
    .config_7_read(config_7_read),
    .config_7_write(config_7_write),
    .config_8_config_addr(config_8_config_addr),
    .config_8_config_data(config_8_config_data),
    .config_8_read(config_8_read),
    .config_8_write(config_8_write),
    .config_9_config_addr(config_9_config_addr),
    .config_9_config_data(config_9_config_data),
    .config_9_read(config_9_read),
    .config_9_write(config_9_write),
    .glb2io_16_X00_Y00(glb2io_16_X00_Y00),
    .glb2io_16_X01_Y00(glb2io_16_X01_Y00),
    .glb2io_16_X02_Y00(glb2io_16_X02_Y00),
    .glb2io_16_X03_Y00(glb2io_16_X03_Y00),
    .glb2io_16_X04_Y00(glb2io_16_X04_Y00),
    .glb2io_16_X05_Y00(glb2io_16_X05_Y00),
    .glb2io_16_X06_Y00(glb2io_16_X06_Y00),
    .glb2io_16_X07_Y00(glb2io_16_X07_Y00),
    .glb2io_16_X08_Y00(glb2io_16_X08_Y00),
    .glb2io_16_X09_Y00(glb2io_16_X09_Y00),
    .glb2io_16_X0A_Y00(glb2io_16_X0A_Y00),
    .glb2io_16_X0B_Y00(glb2io_16_X0B_Y00),
    .glb2io_16_X0C_Y00(glb2io_16_X0C_Y00),
    .glb2io_16_X0D_Y00(glb2io_16_X0D_Y00),
    .glb2io_16_X0E_Y00(glb2io_16_X0E_Y00),
    .glb2io_16_X0F_Y00(glb2io_16_X0F_Y00),
    .glb2io_1_X00_Y00(glb2io_1_X00_Y00),
    .glb2io_1_X01_Y00(glb2io_1_X01_Y00),
    .glb2io_1_X02_Y00(glb2io_1_X02_Y00),
    .glb2io_1_X03_Y00(glb2io_1_X03_Y00),
    .glb2io_1_X04_Y00(glb2io_1_X04_Y00),
    .glb2io_1_X05_Y00(glb2io_1_X05_Y00),
    .glb2io_1_X06_Y00(glb2io_1_X06_Y00),
    .glb2io_1_X07_Y00(glb2io_1_X07_Y00),
    .glb2io_1_X08_Y00(glb2io_1_X08_Y00),
    .glb2io_1_X09_Y00(glb2io_1_X09_Y00),
    .glb2io_1_X0A_Y00(glb2io_1_X0A_Y00),
    .glb2io_1_X0B_Y00(glb2io_1_X0B_Y00),
    .glb2io_1_X0C_Y00(glb2io_1_X0C_Y00),
    .glb2io_1_X0D_Y00(glb2io_1_X0D_Y00),
    .glb2io_1_X0E_Y00(glb2io_1_X0E_Y00),
    .glb2io_1_X0F_Y00(glb2io_1_X0F_Y00),
    .io2glb_16_X00_Y00(Interconnect_inst0_io2glb_16_X00_Y00),
    .io2glb_16_X01_Y00(Interconnect_inst0_io2glb_16_X01_Y00),
    .io2glb_16_X02_Y00(Interconnect_inst0_io2glb_16_X02_Y00),
    .io2glb_16_X03_Y00(Interconnect_inst0_io2glb_16_X03_Y00),
    .io2glb_16_X04_Y00(Interconnect_inst0_io2glb_16_X04_Y00),
    .io2glb_16_X05_Y00(Interconnect_inst0_io2glb_16_X05_Y00),
    .io2glb_16_X06_Y00(Interconnect_inst0_io2glb_16_X06_Y00),
    .io2glb_16_X07_Y00(Interconnect_inst0_io2glb_16_X07_Y00),
    .io2glb_16_X08_Y00(Interconnect_inst0_io2glb_16_X08_Y00),
    .io2glb_16_X09_Y00(Interconnect_inst0_io2glb_16_X09_Y00),
    .io2glb_16_X0A_Y00(Interconnect_inst0_io2glb_16_X0A_Y00),
    .io2glb_16_X0B_Y00(Interconnect_inst0_io2glb_16_X0B_Y00),
    .io2glb_16_X0C_Y00(Interconnect_inst0_io2glb_16_X0C_Y00),
    .io2glb_16_X0D_Y00(Interconnect_inst0_io2glb_16_X0D_Y00),
    .io2glb_16_X0E_Y00(Interconnect_inst0_io2glb_16_X0E_Y00),
    .io2glb_16_X0F_Y00(Interconnect_inst0_io2glb_16_X0F_Y00),
    .io2glb_1_X00_Y00(Interconnect_inst0_io2glb_1_X00_Y00),
    .io2glb_1_X01_Y00(Interconnect_inst0_io2glb_1_X01_Y00),
    .io2glb_1_X02_Y00(Interconnect_inst0_io2glb_1_X02_Y00),
    .io2glb_1_X03_Y00(Interconnect_inst0_io2glb_1_X03_Y00),
    .io2glb_1_X04_Y00(Interconnect_inst0_io2glb_1_X04_Y00),
    .io2glb_1_X05_Y00(Interconnect_inst0_io2glb_1_X05_Y00),
    .io2glb_1_X06_Y00(Interconnect_inst0_io2glb_1_X06_Y00),
    .io2glb_1_X07_Y00(Interconnect_inst0_io2glb_1_X07_Y00),
    .io2glb_1_X08_Y00(Interconnect_inst0_io2glb_1_X08_Y00),
    .io2glb_1_X09_Y00(Interconnect_inst0_io2glb_1_X09_Y00),
    .io2glb_1_X0A_Y00(Interconnect_inst0_io2glb_1_X0A_Y00),
    .io2glb_1_X0B_Y00(Interconnect_inst0_io2glb_1_X0B_Y00),
    .io2glb_1_X0C_Y00(Interconnect_inst0_io2glb_1_X0C_Y00),
    .io2glb_1_X0D_Y00(Interconnect_inst0_io2glb_1_X0D_Y00),
    .io2glb_1_X0E_Y00(Interconnect_inst0_io2glb_1_X0E_Y00),
    .io2glb_1_X0F_Y00(Interconnect_inst0_io2glb_1_X0F_Y00),
    .read_config_data(Interconnect_inst0_read_config_data),
    .reset(reset),
    .stall(stall)
);
assign io2glb_16_X00_Y00 = Interconnect_inst0_io2glb_16_X00_Y00;
assign io2glb_16_X01_Y00 = Interconnect_inst0_io2glb_16_X01_Y00;
assign io2glb_16_X02_Y00 = Interconnect_inst0_io2glb_16_X02_Y00;
assign io2glb_16_X03_Y00 = Interconnect_inst0_io2glb_16_X03_Y00;
assign io2glb_16_X04_Y00 = Interconnect_inst0_io2glb_16_X04_Y00;
assign io2glb_16_X05_Y00 = Interconnect_inst0_io2glb_16_X05_Y00;
assign io2glb_16_X06_Y00 = Interconnect_inst0_io2glb_16_X06_Y00;
assign io2glb_16_X07_Y00 = Interconnect_inst0_io2glb_16_X07_Y00;
assign io2glb_16_X08_Y00 = Interconnect_inst0_io2glb_16_X08_Y00;
assign io2glb_16_X09_Y00 = Interconnect_inst0_io2glb_16_X09_Y00;
assign io2glb_16_X0A_Y00 = Interconnect_inst0_io2glb_16_X0A_Y00;
assign io2glb_16_X0B_Y00 = Interconnect_inst0_io2glb_16_X0B_Y00;
assign io2glb_16_X0C_Y00 = Interconnect_inst0_io2glb_16_X0C_Y00;
assign io2glb_16_X0D_Y00 = Interconnect_inst0_io2glb_16_X0D_Y00;
assign io2glb_16_X0E_Y00 = Interconnect_inst0_io2glb_16_X0E_Y00;
assign io2glb_16_X0F_Y00 = Interconnect_inst0_io2glb_16_X0F_Y00;
assign io2glb_1_X00_Y00 = Interconnect_inst0_io2glb_1_X00_Y00;
assign io2glb_1_X01_Y00 = Interconnect_inst0_io2glb_1_X01_Y00;
assign io2glb_1_X02_Y00 = Interconnect_inst0_io2glb_1_X02_Y00;
assign io2glb_1_X03_Y00 = Interconnect_inst0_io2glb_1_X03_Y00;
assign io2glb_1_X04_Y00 = Interconnect_inst0_io2glb_1_X04_Y00;
assign io2glb_1_X05_Y00 = Interconnect_inst0_io2glb_1_X05_Y00;
assign io2glb_1_X06_Y00 = Interconnect_inst0_io2glb_1_X06_Y00;
assign io2glb_1_X07_Y00 = Interconnect_inst0_io2glb_1_X07_Y00;
assign io2glb_1_X08_Y00 = Interconnect_inst0_io2glb_1_X08_Y00;
assign io2glb_1_X09_Y00 = Interconnect_inst0_io2glb_1_X09_Y00;
assign io2glb_1_X0A_Y00 = Interconnect_inst0_io2glb_1_X0A_Y00;
assign io2glb_1_X0B_Y00 = Interconnect_inst0_io2glb_1_X0B_Y00;
assign io2glb_1_X0C_Y00 = Interconnect_inst0_io2glb_1_X0C_Y00;
assign io2glb_1_X0D_Y00 = Interconnect_inst0_io2glb_1_X0D_Y00;
assign io2glb_1_X0E_Y00 = Interconnect_inst0_io2glb_1_X0E_Y00;
assign io2glb_1_X0F_Y00 = Interconnect_inst0_io2glb_1_X0F_Y00;
assign read_config_data = Interconnect_inst0_read_config_data;
endmodule

