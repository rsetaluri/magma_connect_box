
module Interconnect (
   input  clk,
   output [31:0] read_config_data,
   input  reset,
   input [11:0] stall,

   input [31:0] config_0_config_addr,
   input [31:0] config_0_config_data,
   input [0:0] config_0_read,
   input [0:0] config_0_write,
   input [31:0] config_1_config_addr,
   input [31:0] config_1_config_data,
   input [0:0] config_1_read,
   input [0:0] config_1_write,
   input [31:0] config_2_config_addr,
   input [31:0] config_2_config_data,
   input [0:0] config_2_read,
   input [0:0] config_2_write,
   input [31:0] config_3_config_addr,
   input [31:0] config_3_config_data,
   input [0:0] config_3_read,
   input [0:0] config_3_write,
   input [31:0] config_4_config_addr,
   input [31:0] config_4_config_data,
   input [0:0] config_4_read,
   input [0:0] config_4_write,
   input [31:0] config_5_config_addr,
   input [31:0] config_5_config_data,
   input [0:0] config_5_read,
   input [0:0] config_5_write,
   input [31:0] config_6_config_addr,
   input [31:0] config_6_config_data,
   input [0:0] config_6_read,
   input [0:0] config_6_write,
   input [31:0] config_7_config_addr,
   input [31:0] config_7_config_data,
   input [0:0] config_7_read,
   input [0:0] config_7_write,
   input [31:0] config_8_config_addr,
   input [31:0] config_8_config_data,
   input [0:0] config_8_read,
   input [0:0] config_8_write,
   input [31:0] config_9_config_addr,
   input [31:0] config_9_config_data,
   input [0:0] config_9_read,
   input [0:0] config_9_write,
   input [31:0] config_10_config_addr,
   input [31:0] config_10_config_data,
   input [0:0] config_10_read,
   input [0:0] config_10_write,
   input [31:0] config_11_config_addr,
   input [31:0] config_11_config_data,
   input [0:0] config_11_read,
   input [0:0] config_11_write,
   input [0:0] glb2io_1_X00_Y00,
   output [0:0] io2glb_1_X00_Y00,
   input [15:0] glb2io_16_X00_Y00,
   output [15:0] io2glb_16_X00_Y00,
   input [0:0] glb2io_1_X01_Y00,
   output [0:0] io2glb_1_X01_Y00,
   input [15:0] glb2io_16_X01_Y00,
   output [15:0] io2glb_16_X01_Y00,
   input [0:0] glb2io_1_X02_Y00,
   output [0:0] io2glb_1_X02_Y00,
   input [15:0] glb2io_16_X02_Y00,
   output [15:0] io2glb_16_X02_Y00,
   input [0:0] glb2io_1_X03_Y00,
   output [0:0] io2glb_1_X03_Y00,
   input [15:0] glb2io_16_X03_Y00,
   output [15:0] io2glb_16_X03_Y00,
   input [0:0] glb2io_1_X04_Y00,
   output [0:0] io2glb_1_X04_Y00,
   input [15:0] glb2io_16_X04_Y00,
   output [15:0] io2glb_16_X04_Y00,
   input [0:0] glb2io_1_X05_Y00,
   output [0:0] io2glb_1_X05_Y00,
   input [15:0] glb2io_16_X05_Y00,
   output [15:0] io2glb_16_X05_Y00,
   input [0:0] glb2io_1_X06_Y00,
   output [0:0] io2glb_1_X06_Y00,
   input [15:0] glb2io_16_X06_Y00,
   output [15:0] io2glb_16_X06_Y00,
   input [0:0] glb2io_1_X07_Y00,
   output [0:0] io2glb_1_X07_Y00,
   input [15:0] glb2io_16_X07_Y00,
   output [15:0] io2glb_16_X07_Y00,
   input [0:0] glb2io_1_X08_Y00,
   output [0:0] io2glb_1_X08_Y00,
   input [15:0] glb2io_16_X08_Y00,
   output [15:0] io2glb_16_X08_Y00,
   input [0:0] glb2io_1_X09_Y00,
   output [0:0] io2glb_1_X09_Y00,
   input [15:0] glb2io_16_X09_Y00,
   output [15:0] io2glb_16_X09_Y00,
   input [0:0] glb2io_1_X0A_Y00,
   output [0:0] io2glb_1_X0A_Y00,
   input [15:0] glb2io_16_X0A_Y00,
   output [15:0] io2glb_16_X0A_Y00,
   input [0:0] glb2io_1_X0B_Y00,
   output [0:0] io2glb_1_X0B_Y00,
   input [15:0] glb2io_16_X0B_Y00,
   output [15:0] io2glb_16_X0B_Y00
);
endmodule
